-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 0/Unpack 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_0;
architecture structural of mh_unpack_72_bit_fifo_0 is 
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 0/Unpack 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_1;
architecture structural of mh_unpack_72_bit_fifo_1 is 
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_unpacker_ram_0 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_60_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x71_downto_60_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_unpacker_ram_0;
architecture structural of mh_72_bit_unpacker_ram_0 is 
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal slice_47_down_to_36_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal data_mux_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_24_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal clk_net : std_logic;
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal slice_23_down_to_12_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal write_fifo_0_mux_delay_q_net : std_logic;
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_60_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal write_fifo_1_mux_delay_q_net : std_logic;
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_enable_check_q_net : std_logic_vector( 72-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 1-1 downto 0 );
  signal zero_fifo_value_op_net : std_logic_vector( 72-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  x71_downto_60_fifo_0 <= slice_71_down_to_60_y_net;
  x59_downto_48_fifo_0 <= slice_59_down_to_48_y_net;
  x47_downto_36_fifo_0 <= slice_47_down_to_36_y_net;
  x35_downto_24_fifo_0 <= slice_35_down_to_24_y_net;
  x23_downto_12_fifo_0 <= slice_23_down_to_12_y_net;
  x11_downto_0_fifo_0 <= slice_11_down_to_0_y_net;
  x71_downto_60_fifo_1 <= slice_71_down_to_60_y_net_x0;
  x59_downto_48_fifo_1 <= slice_59_down_to_48_y_net_x0;
  x47_downto_36_fifo_1 <= slice_47_down_to_36_y_net_x0;
  x35_downto_24_fifo_1 <= slice_35_down_to_24_y_net_x0;
  x23_downto_12_fifo_1 <= slice_23_down_to_12_y_net_x0;
  x11_downto_0_fifo_1 <= slice_11_down_to_0_y_net_x0;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_0_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_72_bit_fifo_0 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net,
    x59_downto_48 => slice_59_down_to_48_y_net,
    x47_downto_36 => slice_47_down_to_36_y_net,
    x35_downto_24 => slice_35_down_to_24_y_net,
    x23_downto_12 => slice_23_down_to_12_y_net,
    x11_downto_0 => slice_11_down_to_0_y_net
  );
  unpack_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_72_bit_fifo_1 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net_x0,
    x59_downto_48 => slice_59_down_to_48_y_net_x0,
    x47_downto_36 => slice_47_down_to_36_y_net_x0,
    x35_downto_24 => slice_35_down_to_24_y_net_x0,
    x23_downto_12 => slice_23_down_to_12_y_net_x0,
    x11_downto_0 => slice_11_down_to_0_y_net_x0
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_mux_delay_q_net,
    we => write_fifo_0_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => write_fifo_1_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_q_net
  );
  data_enable_check : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_enable_check_q_net
  );
  data_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_mux_delay_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  enable_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay1_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_0_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_enable_check_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_value_delay_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_998091030b 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_0_empty_net,
    d1(0) => x72bit_frame_fifo_1_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  sync_frame_counter : entity xil_defaultlib.sysgen_counter_4497493dc5 
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_fifo_0_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_0_mux_delay_q_net
  );
  write_fifo_1_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_1_mux_delay_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  zero_fifo_value : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_fifo_value_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => last_value_delay_q_net,
    d1 => zero_fifo_value_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 1/Unpack 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_0_x0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_0_x0;
architecture structural of mh_unpack_72_bit_fifo_0_x0 is 
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 1/Unpack 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_1_x0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_1_x0;
architecture structural of mh_unpack_72_bit_fifo_1_x0 is 
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_unpacker_ram_1 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_60_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x71_downto_60_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_unpacker_ram_1;
architecture structural of mh_72_bit_unpacker_ram_1 is 
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal slice_11_down_to_0_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_60_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal data_enable_check_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal zero_fifo_value_op_net : std_logic_vector( 72-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_mux_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal write_fifo_1_mux_delay_q_net : std_logic;
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal write_fifo_0_mux_delay_q_net : std_logic;
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal data_delay_q_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_60_fifo_0 <= slice_71_down_to_60_y_net;
  x59_downto_48_fifo_0 <= slice_59_down_to_48_y_net;
  x47_downto_36_fifo_0 <= slice_47_down_to_36_y_net;
  x35_downto_24_fifo_0 <= slice_35_down_to_24_y_net;
  x23_downto_12_fifo_0 <= slice_23_down_to_12_y_net;
  x11_downto_0_fifo_0 <= slice_11_down_to_0_y_net;
  x71_downto_60_fifo_1 <= slice_71_down_to_60_y_net_x0;
  x59_downto_48_fifo_1 <= slice_59_down_to_48_y_net_x0;
  x47_downto_36_fifo_1 <= slice_47_down_to_36_y_net_x0;
  x35_downto_24_fifo_1 <= slice_35_down_to_24_y_net_x0;
  x23_downto_12_fifo_1 <= slice_23_down_to_12_y_net_x0;
  x11_downto_0_fifo_1 <= slice_11_down_to_0_y_net_x0;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_1_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_72_bit_fifo_0_x0 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net,
    x59_downto_48 => slice_59_down_to_48_y_net,
    x47_downto_36 => slice_47_down_to_36_y_net,
    x35_downto_24 => slice_35_down_to_24_y_net,
    x23_downto_12 => slice_23_down_to_12_y_net,
    x11_downto_0 => slice_11_down_to_0_y_net
  );
  unpack_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_72_bit_fifo_1_x0 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net_x0,
    x59_downto_48 => slice_59_down_to_48_y_net_x0,
    x47_downto_36 => slice_47_down_to_36_y_net_x0,
    x35_downto_24 => slice_35_down_to_24_y_net_x0,
    x23_downto_12 => slice_23_down_to_12_y_net_x0,
    x11_downto_0 => slice_11_down_to_0_y_net_x0
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_mux_delay_q_net,
    we => write_fifo_0_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => write_fifo_1_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_q_net
  );
  data_enable_check : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_enable_check_q_net
  );
  data_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_mux_delay_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  enable_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay1_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_0_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_enable_check_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_value_delay_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_998091030b 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_0_empty_net,
    d1(0) => x72bit_frame_fifo_1_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  sync_frame_counter : entity xil_defaultlib.sysgen_counter_4497493dc5 
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_fifo_0_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_0_mux_delay_q_net
  );
  write_fifo_1_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_1_mux_delay_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  zero_fifo_value : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_fifo_value_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => last_value_delay_q_net,
    d1 => zero_fifo_value_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 2/Unpack 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_0_x1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_0_x1;
architecture structural of mh_unpack_72_bit_fifo_0_x1 is 
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 2/Unpack 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_1_x1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_1_x1;
architecture structural of mh_unpack_72_bit_fifo_1_x1 is 
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_unpacker_ram_2 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_60_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x71_downto_60_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_unpacker_ram_2;
architecture structural of mh_72_bit_unpacker_ram_2 is 
  signal sync_frame_counter_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal zero_fifo_value_op_net : std_logic_vector( 72-1 downto 0 );
  signal slice_47_down_to_36_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal data_mux_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal write_fifo_1_mux_delay_q_net : std_logic;
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal write_fifo_0_mux_delay_q_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal data_enable_check_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
begin
  x71_downto_60_fifo_0 <= slice_71_down_to_60_y_net;
  x59_downto_48_fifo_0 <= slice_59_down_to_48_y_net;
  x47_downto_36_fifo_0 <= slice_47_down_to_36_y_net;
  x35_downto_24_fifo_0 <= slice_35_down_to_24_y_net;
  x23_downto_12_fifo_0 <= slice_23_down_to_12_y_net;
  x11_downto_0_fifo_0 <= slice_11_down_to_0_y_net;
  x71_downto_60_fifo_1 <= slice_71_down_to_60_y_net_x0;
  x59_downto_48_fifo_1 <= slice_59_down_to_48_y_net_x0;
  x47_downto_36_fifo_1 <= slice_47_down_to_36_y_net_x0;
  x35_downto_24_fifo_1 <= slice_35_down_to_24_y_net_x0;
  x23_downto_12_fifo_1 <= slice_23_down_to_12_y_net_x0;
  x11_downto_0_fifo_1 <= slice_11_down_to_0_y_net_x0;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_2_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_72_bit_fifo_0_x1 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net,
    x59_downto_48 => slice_59_down_to_48_y_net,
    x47_downto_36 => slice_47_down_to_36_y_net,
    x35_downto_24 => slice_35_down_to_24_y_net,
    x23_downto_12 => slice_23_down_to_12_y_net,
    x11_downto_0 => slice_11_down_to_0_y_net
  );
  unpack_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_72_bit_fifo_1_x1 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net_x0,
    x59_downto_48 => slice_59_down_to_48_y_net_x0,
    x47_downto_36 => slice_47_down_to_36_y_net_x0,
    x35_downto_24 => slice_35_down_to_24_y_net_x0,
    x23_downto_12 => slice_23_down_to_12_y_net_x0,
    x11_downto_0 => slice_11_down_to_0_y_net_x0
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_mux_delay_q_net,
    we => write_fifo_0_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => write_fifo_1_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_q_net
  );
  data_enable_check : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_enable_check_q_net
  );
  data_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_mux_delay_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  enable_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay1_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_0_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_enable_check_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_value_delay_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_998091030b 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_0_empty_net,
    d1(0) => x72bit_frame_fifo_1_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  sync_frame_counter : entity xil_defaultlib.sysgen_counter_4497493dc5 
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_fifo_0_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_0_mux_delay_q_net
  );
  write_fifo_1_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_1_mux_delay_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  zero_fifo_value : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_fifo_value_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => last_value_delay_q_net,
    d1 => zero_fifo_value_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 3/Unpack 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_0_x2 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_0_x2;
architecture structural of mh_unpack_72_bit_fifo_0_x2 is 
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 3/Unpack 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_1_x2 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_1_x2;
architecture structural of mh_unpack_72_bit_fifo_1_x2 is 
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_unpacker_ram_3 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_60_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x71_downto_60_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_unpacker_ram_3;
architecture structural of mh_72_bit_unpacker_ram_3 is 
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal write_fifo_0_mux_delay_q_net : std_logic;
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal write_fifo_1_mux_delay_q_net : std_logic;
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal data_mux_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal data_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal data_enable_check_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal zero_fifo_value_op_net : std_logic_vector( 72-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  x71_downto_60_fifo_0 <= slice_71_down_to_60_y_net;
  x59_downto_48_fifo_0 <= slice_59_down_to_48_y_net;
  x47_downto_36_fifo_0 <= slice_47_down_to_36_y_net;
  x35_downto_24_fifo_0 <= slice_35_down_to_24_y_net;
  x23_downto_12_fifo_0 <= slice_23_down_to_12_y_net;
  x11_downto_0_fifo_0 <= slice_11_down_to_0_y_net;
  x71_downto_60_fifo_1 <= slice_71_down_to_60_y_net_x0;
  x59_downto_48_fifo_1 <= slice_59_down_to_48_y_net_x0;
  x47_downto_36_fifo_1 <= slice_47_down_to_36_y_net_x0;
  x35_downto_24_fifo_1 <= slice_35_down_to_24_y_net_x0;
  x23_downto_12_fifo_1 <= slice_23_down_to_12_y_net_x0;
  x11_downto_0_fifo_1 <= slice_11_down_to_0_y_net_x0;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_3_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_72_bit_fifo_0_x2 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net,
    x59_downto_48 => slice_59_down_to_48_y_net,
    x47_downto_36 => slice_47_down_to_36_y_net,
    x35_downto_24 => slice_35_down_to_24_y_net,
    x23_downto_12 => slice_23_down_to_12_y_net,
    x11_downto_0 => slice_11_down_to_0_y_net
  );
  unpack_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_72_bit_fifo_1_x2 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net_x0,
    x59_downto_48 => slice_59_down_to_48_y_net_x0,
    x47_downto_36 => slice_47_down_to_36_y_net_x0,
    x35_downto_24 => slice_35_down_to_24_y_net_x0,
    x23_downto_12 => slice_23_down_to_12_y_net_x0,
    x11_downto_0 => slice_11_down_to_0_y_net_x0
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_mux_delay_q_net,
    we => write_fifo_0_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => write_fifo_1_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_q_net
  );
  data_enable_check : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_enable_check_q_net
  );
  data_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_mux_delay_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  enable_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay1_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_0_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_enable_check_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_value_delay_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_998091030b 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_0_empty_net,
    d1(0) => x72bit_frame_fifo_1_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  sync_frame_counter : entity xil_defaultlib.sysgen_counter_4497493dc5 
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_fifo_0_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_0_mux_delay_q_net
  );
  write_fifo_1_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_1_mux_delay_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  zero_fifo_value : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_fifo_value_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => last_value_delay_q_net,
    d1 => zero_fifo_value_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 4/Unpack 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_0_x3 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_0_x3;
architecture structural of mh_unpack_72_bit_fifo_0_x3 is 
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 4/Unpack 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_72_bit_fifo_1_x3 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_60 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_unpack_72_bit_fifo_1_x3;
architecture structural of mh_unpack_72_bit_fifo_1_x3 is 
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_60 <= slice_71_down_to_60_y_net;
  x59_downto_48 <= slice_59_down_to_48_y_net;
  x47_downto_36 <= slice_47_down_to_36_y_net;
  x35_downto_24 <= slice_35_down_to_24_y_net;
  x23_downto_12 <= slice_23_down_to_12_y_net;
  x11_downto_0 <= slice_11_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_11_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 11,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_11_down_to_0_y_net
  );
  slice_23_down_to_12 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 12,
    new_msb => 23,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_23_down_to_12_y_net
  );
  slice_35_down_to_24 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 24,
    new_msb => 35,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_24_y_net
  );
  slice_47_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 47,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_47_down_to_36_y_net
  );
  slice_59_down_to_48 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 59,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_59_down_to_48_y_net
  );
  slice_71_down_to_60 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 60,
    new_msb => 71,
    x_width => 72,
    y_width => 12
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_60_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/72 Bit Unpacker RAM 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_unpacker_ram_4 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_60_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_0 : out std_logic_vector( 12-1 downto 0 );
    x71_downto_60_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x59_downto_48_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x47_downto_36_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x35_downto_24_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x23_downto_12_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    x11_downto_0_fifo_1 : out std_logic_vector( 12-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_unpacker_ram_4;
architecture structural of mh_72_bit_unpacker_ram_4 is 
  signal data_enable_check_q_net : std_logic_vector( 72-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_23_down_to_12_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal data_in_delay_1_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_60_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal data_mux_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal write_fifo_0_mux_delay_q_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal write_fifo_1_mux_delay_q_net : std_logic;
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_point_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal zero_fifo_value_op_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_60_fifo_0 <= slice_71_down_to_60_y_net;
  x59_downto_48_fifo_0 <= slice_59_down_to_48_y_net;
  x47_downto_36_fifo_0 <= slice_47_down_to_36_y_net;
  x35_downto_24_fifo_0 <= slice_35_down_to_24_y_net;
  x23_downto_12_fifo_0 <= slice_23_down_to_12_y_net;
  x11_downto_0_fifo_0 <= slice_11_down_to_0_y_net;
  x71_downto_60_fifo_1 <= slice_71_down_to_60_y_net_x0;
  x59_downto_48_fifo_1 <= slice_59_down_to_48_y_net_x0;
  x47_downto_36_fifo_1 <= slice_47_down_to_36_y_net_x0;
  x35_downto_24_fifo_1 <= slice_35_down_to_24_y_net_x0;
  x23_downto_12_fifo_1 <= slice_23_down_to_12_y_net_x0;
  x11_downto_0_fifo_1 <= slice_11_down_to_0_y_net_x0;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_4_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_72_bit_fifo_0_x3 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net,
    x59_downto_48 => slice_59_down_to_48_y_net,
    x47_downto_36 => slice_47_down_to_36_y_net,
    x35_downto_24 => slice_35_down_to_24_y_net,
    x23_downto_12 => slice_23_down_to_12_y_net,
    x11_downto_0 => slice_11_down_to_0_y_net
  );
  unpack_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_72_bit_fifo_1_x3 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_60 => slice_71_down_to_60_y_net_x0,
    x59_downto_48 => slice_59_down_to_48_y_net_x0,
    x47_downto_36 => slice_47_down_to_36_y_net_x0,
    x35_downto_24 => slice_35_down_to_24_y_net_x0,
    x23_downto_12 => slice_23_down_to_12_y_net_x0,
    x11_downto_0 => slice_11_down_to_0_y_net_x0
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_mux_delay_q_net,
    we => write_fifo_0_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => write_fifo_1_mux_delay_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_point_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_q_net
  );
  data_enable_check : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_enable_check_q_net
  );
  data_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_mux_delay_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  last_point_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => last_point_delay_1_q_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_0_op_net,
    d1 => last_point_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => last_point_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_enable_check_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_value_delay_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_998091030b 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_0_empty_net,
    d1(0) => x72bit_frame_fifo_1_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_6a55809cad 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  sync_frame_counter : entity xil_defaultlib.sysgen_counter_4497493dc5 
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_fifo_0_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_0_mux_delay_q_net
  );
  write_fifo_1_mux_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => write_fifo_1_mux_delay_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  zero_fifo_value : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_fifo_value_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => last_value_delay_q_net,
    d1 => zero_fifo_value_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer/Data Point Tracker
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_data_point_tracker is
  port (
    data_in_ram_0 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_1 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_2 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_3 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_4 : in std_logic_vector( 72-1 downto 0 );
    valid_enable_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_out_ram_0 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_1 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_2 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_3 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_4 : out std_logic_vector( 72-1 downto 0 );
    valid_enable_out : out std_logic_vector( 1-1 downto 0 );
    last_value_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_data_point_tracker;
architecture structural of mh_data_point_tracker is 
  signal valid_delay_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_point_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_data_point_value_op_net : std_logic_vector( 7-1 downto 0 );
  signal data_point_counter_op_net : std_logic_vector( 7-1 downto 0 );
  signal data_in_delay_1_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal clk_net : std_logic;
  signal data_in_delay_0_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_0_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_0_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_0_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_0_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
begin
  data_out_ram_0 <= data_in_delay_1_ram_0_q_net;
  data_out_ram_1 <= data_in_delay_1_ram_1_q_net;
  data_out_ram_2 <= data_in_delay_1_ram_2_q_net;
  data_out_ram_3 <= data_in_delay_1_ram_3_q_net;
  data_out_ram_4 <= data_in_delay_1_ram_4_q_net;
  valid_enable_out <= valid_delay_1_q_net;
  last_value_out <= last_value_enable_y_net;
  dual_port_ram_0_douta_net <= data_in_ram_0;
  dual_port_ram_1_douta_net <= data_in_ram_1;
  dual_port_ram_2_douta_net <= data_in_ram_2;
  dual_port_ram_3_douta_net <= data_in_ram_3;
  dual_port_ram_4_douta_net <= data_in_ram_4;
  convert_to_bool_dout_net <= valid_enable_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  data_in_delay_0_ram_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_0_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_0_q_net
  );
  data_in_delay_0_ram_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_1_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_1_q_net
  );
  data_in_delay_0_ram_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_2_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_2_q_net
  );
  data_in_delay_0_ram_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_3_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_3_q_net
  );
  data_in_delay_0_ram_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_4_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_4_q_net
  );
  data_in_delay_1_ram_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_0_q_net
  );
  data_in_delay_1_ram_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_1_q_net
  );
  data_in_delay_1_ram_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_2_q_net
  );
  data_in_delay_1_ram_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_3_q_net
  );
  data_in_delay_1_ram_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_4_q_net
  );
  data_point_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 66,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i0",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    rst => "0",
    clr => '0',
    en => convert_to_bool_dout_net,
    clk => clk_net,
    ce => ce_net,
    op => data_point_counter_op_net
  );
  last_data_point_value : entity xil_defaultlib.sysgen_constant_6b755964f8 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => last_data_point_value_op_net
  );
  last_point : entity xil_defaultlib.sysgen_relational_d18eb5aea1 
  port map (
    clr => '0',
    a => data_point_counter_op_net,
    b => last_data_point_value_op_net,
    clk => clk_net,
    ce => ce_net,
    op => last_point_op_net
  );
  last_value_enable : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => valid_delay_0_q_net,
    d1 => last_point_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_enable_y_net
  );
  valid_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_to_bool_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_delay_0_q_net
  );
  valid_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_delay_1_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Frame RAM Slicer
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_frame_ram_slicer is
  port (
    data_in_ram_0 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_1 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_2 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_3 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_4 : in std_logic_vector( 72-1 downto 0 );
    valid_in : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    frame_12_bit_bin_value_0_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11_ram_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_0_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11_ram_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_0_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11_ram_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_0_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11_ram_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_0_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10_ram_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11_ram_4 : out std_logic_vector( 12-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_0 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_1 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_2 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_3 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_4 : out std_logic_vector( 1-1 downto 0 )
  );
end mh_frame_ram_slicer;
architecture structural of mh_frame_ram_slicer is 
  signal delay_47_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_60_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_47_down_to_36_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net : std_logic_vector( 12-1 downto 0 );
  signal data_in_delay_1_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_59_down_to_48_y_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 12-1 downto 0 );
  signal valid_sync_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_11_down_to_0_y_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal data_in_delay_1_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal valid_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal slice_59_down_to_48_y_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal slice_11_down_to_0_y_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice_35_down_to_24_y_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal slice_71_down_to_60_y_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal data_in_delay_1_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_24_y_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal slice_35_down_to_24_y_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal slice_23_down_to_12_y_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal valid_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal slice_11_down_to_0_y_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal data_in_delay_1_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_60_y_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal slice_59_down_to_48_y_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal slice_47_down_to_36_y_net_x6 : std_logic_vector( 12-1 downto 0 );
begin
  frame_12_bit_bin_value_0_ram_0 <= delay_5_q_net;
  frame_12_bit_bin_value_1_ram_0 <= delay_4_q_net;
  frame_12_bit_bin_value_2_ram_0 <= delay_3_q_net;
  frame_12_bit_bin_value_3_ram_0 <= delay_2_q_net;
  frame_12_bit_bin_value_4_ram_0 <= delay_1_q_net;
  frame_12_bit_bin_value_5_ram_0 <= delay_0_q_net;
  frame_12_bit_bin_value_6_ram_0 <= delay_11_q_net;
  frame_12_bit_bin_value_7_ram_0 <= delay_10_q_net;
  frame_12_bit_bin_value_8_ram_0 <= delay_9_q_net;
  frame_12_bit_bin_value_9_ram_0 <= delay_8_q_net;
  frame_12_bit_bin_value_10_ram_0 <= delay_7_q_net;
  frame_12_bit_bin_value_11_ram_0 <= delay_6_q_net;
  frame_12_bit_bin_value_0_ram_1 <= delay_19_q_net;
  frame_12_bit_bin_value_1_ram_1 <= delay_18_q_net;
  frame_12_bit_bin_value_2_ram_1 <= delay_17_q_net;
  frame_12_bit_bin_value_3_ram_1 <= delay_16_q_net;
  frame_12_bit_bin_value_4_ram_1 <= delay_13_q_net;
  frame_12_bit_bin_value_5_ram_1 <= delay_12_q_net;
  frame_12_bit_bin_value_6_ram_1 <= delay_15_q_net;
  frame_12_bit_bin_value_7_ram_1 <= delay_14_q_net;
  frame_12_bit_bin_value_8_ram_1 <= delay_23_q_net;
  frame_12_bit_bin_value_9_ram_1 <= delay_22_q_net;
  frame_12_bit_bin_value_10_ram_1 <= delay_21_q_net;
  frame_12_bit_bin_value_11_ram_1 <= delay_20_q_net;
  frame_12_bit_bin_value_0_ram_2 <= delay_43_q_net;
  frame_12_bit_bin_value_1_ram_2 <= delay_42_q_net;
  frame_12_bit_bin_value_2_ram_2 <= delay_41_q_net;
  frame_12_bit_bin_value_3_ram_2 <= delay_36_q_net;
  frame_12_bit_bin_value_4_ram_2 <= delay_25_q_net;
  frame_12_bit_bin_value_5_ram_2 <= delay_24_q_net;
  frame_12_bit_bin_value_6_ram_2 <= delay_27_q_net;
  frame_12_bit_bin_value_7_ram_2 <= delay_26_q_net;
  frame_12_bit_bin_value_8_ram_2 <= delay_47_q_net;
  frame_12_bit_bin_value_9_ram_2 <= delay_46_q_net;
  frame_12_bit_bin_value_10_ram_2 <= delay_45_q_net;
  frame_12_bit_bin_value_11_ram_2 <= delay_44_q_net;
  frame_12_bit_bin_value_0_ram_3 <= delay_35_q_net;
  frame_12_bit_bin_value_1_ram_3 <= delay_34_q_net;
  frame_12_bit_bin_value_2_ram_3 <= delay_33_q_net;
  frame_12_bit_bin_value_3_ram_3 <= delay_32_q_net;
  frame_12_bit_bin_value_4_ram_3 <= delay_29_q_net;
  frame_12_bit_bin_value_5_ram_3 <= delay_28_q_net;
  frame_12_bit_bin_value_6_ram_3 <= delay_31_q_net;
  frame_12_bit_bin_value_7_ram_3 <= delay_30_q_net;
  frame_12_bit_bin_value_8_ram_3 <= delay_40_q_net;
  frame_12_bit_bin_value_9_ram_3 <= delay_39_q_net;
  frame_12_bit_bin_value_10_ram_3 <= delay_38_q_net;
  frame_12_bit_bin_value_11_ram_3 <= delay_37_q_net;
  frame_12_bit_bin_value_0_ram_4 <= delay_67_q_net;
  frame_12_bit_bin_value_1_ram_4 <= delay_66_q_net;
  frame_12_bit_bin_value_2_ram_4 <= delay_65_q_net;
  frame_12_bit_bin_value_3_ram_4 <= delay_60_q_net;
  frame_12_bit_bin_value_4_ram_4 <= delay_49_q_net;
  frame_12_bit_bin_value_5_ram_4 <= delay_48_q_net;
  frame_12_bit_bin_value_6_ram_4 <= delay_51_q_net;
  frame_12_bit_bin_value_7_ram_4 <= delay_50_q_net;
  frame_12_bit_bin_value_8_ram_4 <= delay_71_q_net;
  frame_12_bit_bin_value_9_ram_4 <= delay_70_q_net;
  frame_12_bit_bin_value_10_ram_4 <= delay_69_q_net;
  frame_12_bit_bin_value_11_ram_4 <= delay_68_q_net;
  valid_out <= valid_sync_y_net;
  wrote_to_last_fifo_ram_0 <= logical_y_net_x3;
  wrote_to_last_fifo_ram_1 <= logical_y_net_x2;
  wrote_to_last_fifo_ram_2 <= logical_y_net_x1;
  wrote_to_last_fifo_ram_3 <= logical_y_net_x0;
  wrote_to_last_fifo_ram_4 <= logical_y_net;
  dual_port_ram_0_douta_net <= data_in_ram_0;
  dual_port_ram_1_douta_net <= data_in_ram_1;
  dual_port_ram_2_douta_net <= data_in_ram_2;
  dual_port_ram_3_douta_net <= data_in_ram_3;
  dual_port_ram_4_douta_net <= data_in_ram_4;
  convert_to_bool_dout_net <= valid_in;
  read_out_y_net <= read_enable;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x72_bit_unpacker_ram_0 : entity xil_defaultlib.mh_72_bit_unpacker_ram_0 
  port map (
    data_in => data_in_delay_1_ram_0_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_60_fifo_0 => slice_71_down_to_60_y_net_x8,
    x59_downto_48_fifo_0 => slice_59_down_to_48_y_net_x8,
    x47_downto_36_fifo_0 => slice_47_down_to_36_y_net_x8,
    x35_downto_24_fifo_0 => slice_35_down_to_24_y_net_x8,
    x23_downto_12_fifo_0 => slice_23_down_to_12_y_net_x8,
    x11_downto_0_fifo_0 => slice_11_down_to_0_y_net_x8,
    x71_downto_60_fifo_1 => slice_71_down_to_60_y_net_x7,
    x59_downto_48_fifo_1 => slice_59_down_to_48_y_net_x7,
    x47_downto_36_fifo_1 => slice_47_down_to_36_y_net_x7,
    x35_downto_24_fifo_1 => slice_35_down_to_24_y_net_x7,
    x23_downto_12_fifo_1 => slice_23_down_to_12_y_net_x7,
    x11_downto_0_fifo_1 => slice_11_down_to_0_y_net_x7,
    valid_out => valid_q_net_x3,
    wrote_to_a_fifo => logical_y_net_x3
  );
  x72_bit_unpacker_ram_1 : entity xil_defaultlib.mh_72_bit_unpacker_ram_1 
  port map (
    data_in => data_in_delay_1_ram_1_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_60_fifo_0 => slice_71_down_to_60_y_net_x6,
    x59_downto_48_fifo_0 => slice_59_down_to_48_y_net_x6,
    x47_downto_36_fifo_0 => slice_47_down_to_36_y_net_x6,
    x35_downto_24_fifo_0 => slice_35_down_to_24_y_net_x6,
    x23_downto_12_fifo_0 => slice_23_down_to_12_y_net_x6,
    x11_downto_0_fifo_0 => slice_11_down_to_0_y_net_x6,
    x71_downto_60_fifo_1 => slice_71_down_to_60_y_net_x5,
    x59_downto_48_fifo_1 => slice_59_down_to_48_y_net_x5,
    x47_downto_36_fifo_1 => slice_47_down_to_36_y_net_x5,
    x35_downto_24_fifo_1 => slice_35_down_to_24_y_net_x5,
    x23_downto_12_fifo_1 => slice_23_down_to_12_y_net_x5,
    x11_downto_0_fifo_1 => slice_11_down_to_0_y_net_x5,
    valid_out => valid_q_net_x2,
    wrote_to_a_fifo => logical_y_net_x2
  );
  x72_bit_unpacker_ram_2 : entity xil_defaultlib.mh_72_bit_unpacker_ram_2 
  port map (
    data_in => data_in_delay_1_ram_2_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_60_fifo_0 => slice_71_down_to_60_y_net_x4,
    x59_downto_48_fifo_0 => slice_59_down_to_48_y_net_x4,
    x47_downto_36_fifo_0 => slice_47_down_to_36_y_net_x4,
    x35_downto_24_fifo_0 => slice_35_down_to_24_y_net_x4,
    x23_downto_12_fifo_0 => slice_23_down_to_12_y_net_x4,
    x11_downto_0_fifo_0 => slice_11_down_to_0_y_net_x4,
    x71_downto_60_fifo_1 => slice_71_down_to_60_y_net_x3,
    x59_downto_48_fifo_1 => slice_59_down_to_48_y_net_x3,
    x47_downto_36_fifo_1 => slice_47_down_to_36_y_net_x3,
    x35_downto_24_fifo_1 => slice_35_down_to_24_y_net_x3,
    x23_downto_12_fifo_1 => slice_23_down_to_12_y_net_x3,
    x11_downto_0_fifo_1 => slice_11_down_to_0_y_net_x3,
    valid_out => valid_q_net_x1,
    wrote_to_a_fifo => logical_y_net_x1
  );
  x72_bit_unpacker_ram_3 : entity xil_defaultlib.mh_72_bit_unpacker_ram_3 
  port map (
    data_in => data_in_delay_1_ram_3_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_60_fifo_0 => slice_71_down_to_60_y_net_x2,
    x59_downto_48_fifo_0 => slice_59_down_to_48_y_net_x2,
    x47_downto_36_fifo_0 => slice_47_down_to_36_y_net_x2,
    x35_downto_24_fifo_0 => slice_35_down_to_24_y_net_x2,
    x23_downto_12_fifo_0 => slice_23_down_to_12_y_net_x2,
    x11_downto_0_fifo_0 => slice_11_down_to_0_y_net_x2,
    x71_downto_60_fifo_1 => slice_71_down_to_60_y_net_x1,
    x59_downto_48_fifo_1 => slice_59_down_to_48_y_net_x1,
    x47_downto_36_fifo_1 => slice_47_down_to_36_y_net_x1,
    x35_downto_24_fifo_1 => slice_35_down_to_24_y_net_x1,
    x23_downto_12_fifo_1 => slice_23_down_to_12_y_net_x1,
    x11_downto_0_fifo_1 => slice_11_down_to_0_y_net_x1,
    valid_out => valid_q_net_x0,
    wrote_to_a_fifo => logical_y_net_x0
  );
  x72_bit_unpacker_ram_4 : entity xil_defaultlib.mh_72_bit_unpacker_ram_4 
  port map (
    data_in => data_in_delay_1_ram_4_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_60_fifo_0 => slice_71_down_to_60_y_net_x0,
    x59_downto_48_fifo_0 => slice_59_down_to_48_y_net_x0,
    x47_downto_36_fifo_0 => slice_47_down_to_36_y_net_x0,
    x35_downto_24_fifo_0 => slice_35_down_to_24_y_net_x0,
    x23_downto_12_fifo_0 => slice_23_down_to_12_y_net_x0,
    x11_downto_0_fifo_0 => slice_11_down_to_0_y_net_x0,
    x71_downto_60_fifo_1 => slice_71_down_to_60_y_net,
    x59_downto_48_fifo_1 => slice_59_down_to_48_y_net,
    x47_downto_36_fifo_1 => slice_47_down_to_36_y_net,
    x35_downto_24_fifo_1 => slice_35_down_to_24_y_net,
    x23_downto_12_fifo_1 => slice_23_down_to_12_y_net,
    x11_downto_0_fifo_1 => slice_11_down_to_0_y_net,
    valid_out => valid_q_net,
    wrote_to_a_fifo => logical_y_net
  );
  data_point_tracker : entity xil_defaultlib.mh_data_point_tracker 
  port map (
    data_in_ram_0 => dual_port_ram_0_douta_net,
    data_in_ram_1 => dual_port_ram_1_douta_net,
    data_in_ram_2 => dual_port_ram_2_douta_net,
    data_in_ram_3 => dual_port_ram_3_douta_net,
    data_in_ram_4 => dual_port_ram_4_douta_net,
    valid_enable_in => convert_to_bool_dout_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    data_out_ram_0 => data_in_delay_1_ram_0_q_net,
    data_out_ram_1 => data_in_delay_1_ram_1_q_net,
    data_out_ram_2 => data_in_delay_1_ram_2_q_net,
    data_out_ram_3 => data_in_delay_1_ram_3_q_net,
    data_out_ram_4 => data_in_delay_1_ram_4_q_net,
    valid_enable_out => valid_delay_1_q_net,
    last_value_out => last_value_enable_y_net
  );
  delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_0_q_net
  );
  delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_1_q_net
  );
  delay_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_10_q_net
  );
  delay_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_11_q_net
  );
  delay_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_12_q_net
  );
  delay_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_13_q_net
  );
  delay_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_14_q_net
  );
  delay_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_15_q_net
  );
  delay_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_16_q_net
  );
  delay_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_17_q_net
  );
  delay_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_18_q_net
  );
  delay_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_19_q_net
  );
  delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_2_q_net
  );
  delay_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_20_q_net
  );
  delay_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_21_q_net
  );
  delay_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_22_q_net
  );
  delay_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_23_q_net
  );
  delay_24 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_24_q_net
  );
  delay_25 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_25_q_net
  );
  delay_26 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_26_q_net
  );
  delay_27 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_27_q_net
  );
  delay_28 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_28_q_net
  );
  delay_29 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_29_q_net
  );
  delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_3_q_net
  );
  delay_30 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_30_q_net
  );
  delay_31 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_31_q_net
  );
  delay_32 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_32_q_net
  );
  delay_33 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_33_q_net
  );
  delay_34 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_34_q_net
  );
  delay_35 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_35_q_net
  );
  delay_36 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_36_q_net
  );
  delay_37 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_37_q_net
  );
  delay_38 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_38_q_net
  );
  delay_39 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_39_q_net
  );
  delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_4_q_net
  );
  delay_40 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_40_q_net
  );
  delay_41 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_41_q_net
  );
  delay_42 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_42_q_net
  );
  delay_43 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_43_q_net
  );
  delay_44 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_44_q_net
  );
  delay_45 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_45_q_net
  );
  delay_46 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_46_q_net
  );
  delay_47 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_47_q_net
  );
  delay_48 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_48_q_net
  );
  delay_49 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_49_q_net
  );
  delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_5_q_net
  );
  delay_50 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_50_q_net
  );
  delay_51 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_51_q_net
  );
  delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_6_q_net
  );
  delay_60 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_60_q_net
  );
  delay_65 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_65_q_net
  );
  delay_66 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_23_down_to_12_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_66_q_net
  );
  delay_67 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_11_down_to_0_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_67_q_net
  );
  delay_68 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_60_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_68_q_net
  );
  delay_69 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_69_q_net
  );
  delay_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_59_down_to_48_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_7_q_net
  );
  delay_70 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_70_q_net
  );
  delay_71 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_71_q_net
  );
  delay_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_47_down_to_36_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_8_q_net
  );
  delay_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_24_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_9_q_net
  );
  valid_sync : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => valid_q_net_x3,
    d1 => valid_q_net_x2,
    d2 => valid_q_net_x1,
    d3 => valid_q_net_x0,
    d4 => valid_q_net,
    clk => clk_net,
    ce => ce_net,
    y => valid_sync_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 0/Unpack Kernel 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_0;
architecture structural of mh_unpack_kernel_72_bit_fifo_0 is 
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 0/Unpack Kernel 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_1;
architecture structural of mh_unpack_kernel_72_bit_fifo_1 is 
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 0/Unpack Kernel 72 Bit FIFO 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_2 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_2;
architecture structural of mh_unpack_kernel_72_bit_fifo_2 is 
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_2_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_kernel_unpacker_ram_0 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_54_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_kernel_unpacker_ram_0;
architecture structural of mh_72_bit_kernel_unpacker_ram_0 is 
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_54_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_53_down_to_36_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal last_fifo_written_to_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal clk_net : std_logic;
  signal slice_17_down_to_0_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal slice_53_down_to_36_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal data_delay_4_q_net : std_logic;
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal data_delay_5_q_net : std_logic;
  signal data_delay_6_q_net : std_logic;
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal x72bit_frame_fifo_2_empty_net : std_logic;
  signal x72bit_frame_fifo_2_full_net : std_logic;
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_point_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_2_op_net : std_logic_vector( 2-1 downto 0 );
  signal write_to_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_fifo_written_to_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_7_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 2-1 downto 0 );
  signal zero_out_op_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_54_fifo_0 <= slice_71_down_to_54_y_net;
  x53_downto_36_fifo_0 <= slice_53_down_to_36_y_net;
  x35_downto_18_fifo_0 <= slice_35_down_to_18_y_net;
  x17_downto_0_fifo_0 <= slice_17_down_to_0_y_net;
  x71_downto_54_fifo_1 <= slice_71_down_to_54_y_net_x0;
  x53_downto_36_fifo_1 <= slice_53_down_to_36_y_net_x0;
  x35_downto_18_fifo_1 <= slice_35_down_to_18_y_net_x0;
  x17_downto_0_fifo_1 <= slice_17_down_to_0_y_net_x0;
  x71_downto_54_fifo_2 <= slice_71_down_to_54_y_net_x1;
  x53_downto_36_fifo_2 <= slice_53_down_to_36_y_net_x1;
  x35_downto_18_fifo_2 <= slice_35_down_to_18_y_net_x1;
  x17_downto_0_fifo_2 <= slice_17_down_to_0_y_net_x1;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  wrote_to_last_fifo <= last_fifo_written_to_1_q_net;
  data_in_delay_1_ram_0_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_kernel_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_0 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net,
    x53_downto_36 => slice_53_down_to_36_y_net,
    x35_downto_18 => slice_35_down_to_18_y_net,
    x17_downto_0 => slice_17_down_to_0_y_net
  );
  unpack_kernel_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_1 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x0,
    x53_downto_36 => slice_53_down_to_36_y_net_x0,
    x35_downto_18 => slice_35_down_to_18_y_net_x0,
    x17_downto_0 => slice_17_down_to_0_y_net_x0
  );
  unpack_kernel_72_bit_fifo_2 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_2 
  port map (
    x72_bit_input => x72bit_frame_fifo_2_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x1,
    x53_downto_36 => slice_53_down_to_36_y_net_x1,
    x35_downto_18 => slice_35_down_to_18_y_net_x1,
    x17_downto_0 => slice_17_down_to_0_y_net_x1
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_delay_3_q_net,
    we => data_delay_4_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_5_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  x72bit_frame_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_6_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_2_dout_net,
    empty => x72bit_frame_fifo_2_empty_net,
    full => x72bit_frame_fifo_2_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  data_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_0_q_net
  );
  data_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_1_q_net
  );
  data_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_2_q_net
  );
  data_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_3_q_net
  );
  data_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_4_q_net
  );
  data_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_5_q_net
  );
  data_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_6_q_net
  );
  data_delay_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_7_q_net
  );
  data_delay_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_8_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  fifo_2 : entity xil_defaultlib.sysgen_constant_9d2d62a34e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_2_op_net
  );
  last_fifo_written_to : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d(0) => data_delay_6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_fifo_written_to_q_net
  );
  last_fifo_written_to_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_fifo_written_to_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_fifo_written_to_1_q_net
  );
  last_point_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => last_point_delay_q_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => last_point_delay_q_net,
    d1 => store_in_fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_bypass_fifo_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_2_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_2_y_net
  );
  logical : entity xil_defaultlib.sysgen_logical_17bd555d9a 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_1_empty_net,
    d1(0) => x72bit_frame_fifo_2_empty_net,
    d2(0) => x72bit_frame_fifo_0_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  store_in_fifo_2 : entity xil_defaultlib.sysgen_relational_bf21415019 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_2_op_net
  );
  sync_frame_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  write_to_fifo_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_2_y_net
  );
  zero_out : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_out_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => data_delay_8_q_net,
    d0 => data_delay_2_q_net,
    d1 => zero_out_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 1/Unpack Kernel 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_0_x0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_0_x0;
architecture structural of mh_unpack_kernel_72_bit_fifo_0_x0 is 
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 1/Unpack Kernel 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_1_x0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_1_x0;
architecture structural of mh_unpack_kernel_72_bit_fifo_1_x0 is 
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 1/Unpack Kernel 72 Bit FIFO 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_2_x0 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_2_x0;
architecture structural of mh_unpack_kernel_72_bit_fifo_2_x0 is 
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_2_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_kernel_unpacker_ram_1 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_54_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_kernel_unpacker_ram_1;
architecture structural of mh_72_bit_kernel_unpacker_ram_1 is 
  signal slice_71_down_to_54_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal data_in_delay_1_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_35_down_to_18_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal slice_35_down_to_18_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal data_delay_6_q_net : std_logic;
  signal data_delay_4_q_net : std_logic;
  signal data_delay_5_q_net : std_logic;
  signal x72bit_frame_fifo_2_full_net : std_logic;
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_2_empty_net : std_logic;
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_point_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_2_op_net : std_logic_vector( 2-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 2-1 downto 0 );
  signal store_in_fifo_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal zero_out_op_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_54_fifo_0 <= slice_71_down_to_54_y_net;
  x53_downto_36_fifo_0 <= slice_53_down_to_36_y_net;
  x35_downto_18_fifo_0 <= slice_35_down_to_18_y_net;
  x17_downto_0_fifo_0 <= slice_17_down_to_0_y_net;
  x71_downto_54_fifo_1 <= slice_71_down_to_54_y_net_x0;
  x53_downto_36_fifo_1 <= slice_53_down_to_36_y_net_x0;
  x35_downto_18_fifo_1 <= slice_35_down_to_18_y_net_x0;
  x17_downto_0_fifo_1 <= slice_17_down_to_0_y_net_x0;
  x71_downto_54_fifo_2 <= slice_71_down_to_54_y_net_x1;
  x53_downto_36_fifo_2 <= slice_53_down_to_36_y_net_x1;
  x35_downto_18_fifo_2 <= slice_35_down_to_18_y_net_x1;
  x17_downto_0_fifo_2 <= slice_17_down_to_0_y_net_x1;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_1_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_kernel_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_0_x0 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net,
    x53_downto_36 => slice_53_down_to_36_y_net,
    x35_downto_18 => slice_35_down_to_18_y_net,
    x17_downto_0 => slice_17_down_to_0_y_net
  );
  unpack_kernel_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_1_x0 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x0,
    x53_downto_36 => slice_53_down_to_36_y_net_x0,
    x35_downto_18 => slice_35_down_to_18_y_net_x0,
    x17_downto_0 => slice_17_down_to_0_y_net_x0
  );
  unpack_kernel_72_bit_fifo_2 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_2_x0 
  port map (
    x72_bit_input => x72bit_frame_fifo_2_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x1,
    x53_downto_36 => slice_53_down_to_36_y_net_x1,
    x35_downto_18 => slice_35_down_to_18_y_net_x1,
    x17_downto_0 => slice_17_down_to_0_y_net_x1
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_delay_3_q_net,
    we => data_delay_4_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_5_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  x72bit_frame_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_6_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_2_dout_net,
    empty => x72bit_frame_fifo_2_empty_net,
    full => x72bit_frame_fifo_2_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_0_q_net
  );
  data_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_1_q_net
  );
  data_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_2_q_net
  );
  data_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_3_q_net
  );
  data_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_4_q_net
  );
  data_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_5_q_net
  );
  data_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_6_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  fifo_2 : entity xil_defaultlib.sysgen_constant_9d2d62a34e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_2_op_net
  );
  last_point_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => last_point_delay_q_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => last_point_delay_q_net,
    d1 => store_in_fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_bypass_fifo_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_2_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_2_y_net
  );
  logical : entity xil_defaultlib.sysgen_logical_17bd555d9a 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_1_empty_net,
    d1(0) => x72bit_frame_fifo_2_empty_net,
    d2(0) => x72bit_frame_fifo_0_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  store_in_fifo_2 : entity xil_defaultlib.sysgen_relational_bf21415019 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_2_op_net
  );
  sync_frame_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  write_to_fifo_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_2_y_net
  );
  zero_out : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_out_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => data_delay_2_q_net,
    d1 => zero_out_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 2/Unpack Kernel 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_0_x1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_0_x1;
architecture structural of mh_unpack_kernel_72_bit_fifo_0_x1 is 
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 2/Unpack Kernel 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_1_x1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_1_x1;
architecture structural of mh_unpack_kernel_72_bit_fifo_1_x1 is 
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 2/Unpack Kernel 72 Bit FIFO 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_2_x1 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_2_x1;
architecture structural of mh_unpack_kernel_72_bit_fifo_2_x1 is 
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_2_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_kernel_unpacker_ram_2 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_54_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_kernel_unpacker_ram_2;
architecture structural of mh_72_bit_kernel_unpacker_ram_2 is 
  signal slice_35_down_to_18_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_2_full_net : std_logic;
  signal data_delay_6_q_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal data_delay_4_q_net : std_logic;
  signal ce_net : std_logic;
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal data_delay_5_q_net : std_logic;
  signal x72bit_frame_fifo_2_empty_net : std_logic;
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_point_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_2_op_net : std_logic_vector( 2-1 downto 0 );
  signal last_value_bypass_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 2-1 downto 0 );
  signal zero_out_op_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_54_fifo_0 <= slice_71_down_to_54_y_net;
  x53_downto_36_fifo_0 <= slice_53_down_to_36_y_net;
  x35_downto_18_fifo_0 <= slice_35_down_to_18_y_net;
  x17_downto_0_fifo_0 <= slice_17_down_to_0_y_net;
  x71_downto_54_fifo_1 <= slice_71_down_to_54_y_net_x0;
  x53_downto_36_fifo_1 <= slice_53_down_to_36_y_net_x0;
  x35_downto_18_fifo_1 <= slice_35_down_to_18_y_net_x0;
  x17_downto_0_fifo_1 <= slice_17_down_to_0_y_net_x0;
  x71_downto_54_fifo_2 <= slice_71_down_to_54_y_net_x1;
  x53_downto_36_fifo_2 <= slice_53_down_to_36_y_net_x1;
  x35_downto_18_fifo_2 <= slice_35_down_to_18_y_net_x1;
  x17_downto_0_fifo_2 <= slice_17_down_to_0_y_net_x1;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_2_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_kernel_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_0_x1 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net,
    x53_downto_36 => slice_53_down_to_36_y_net,
    x35_downto_18 => slice_35_down_to_18_y_net,
    x17_downto_0 => slice_17_down_to_0_y_net
  );
  unpack_kernel_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_1_x1 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x0,
    x53_downto_36 => slice_53_down_to_36_y_net_x0,
    x35_downto_18 => slice_35_down_to_18_y_net_x0,
    x17_downto_0 => slice_17_down_to_0_y_net_x0
  );
  unpack_kernel_72_bit_fifo_2 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_2_x1 
  port map (
    x72_bit_input => x72bit_frame_fifo_2_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x1,
    x53_downto_36 => slice_53_down_to_36_y_net_x1,
    x35_downto_18 => slice_35_down_to_18_y_net_x1,
    x17_downto_0 => slice_17_down_to_0_y_net_x1
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_delay_3_q_net,
    we => data_delay_4_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_5_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  x72bit_frame_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_6_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_2_dout_net,
    empty => x72bit_frame_fifo_2_empty_net,
    full => x72bit_frame_fifo_2_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_0_q_net
  );
  data_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_1_q_net
  );
  data_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_2_q_net
  );
  data_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_3_q_net
  );
  data_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_4_q_net
  );
  data_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_5_q_net
  );
  data_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_6_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  fifo_2 : entity xil_defaultlib.sysgen_constant_9d2d62a34e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_2_op_net
  );
  last_point_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => last_point_delay_q_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => last_point_delay_q_net,
    d1 => store_in_fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_bypass_fifo_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_2_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_2_y_net
  );
  logical : entity xil_defaultlib.sysgen_logical_17bd555d9a 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_1_empty_net,
    d1(0) => x72bit_frame_fifo_2_empty_net,
    d2(0) => x72bit_frame_fifo_0_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  store_in_fifo_2 : entity xil_defaultlib.sysgen_relational_bf21415019 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_2_op_net
  );
  sync_frame_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  write_to_fifo_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_2_y_net
  );
  zero_out : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_out_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => data_delay_2_q_net,
    d1 => zero_out_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 3/Unpack Kernel 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_0_x2 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_0_x2;
architecture structural of mh_unpack_kernel_72_bit_fifo_0_x2 is 
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 3/Unpack Kernel 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_1_x2 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_1_x2;
architecture structural of mh_unpack_kernel_72_bit_fifo_1_x2 is 
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 3/Unpack Kernel 72 Bit FIFO 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_2_x2 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_2_x2;
architecture structural of mh_unpack_kernel_72_bit_fifo_2_x2 is 
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_2_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_kernel_unpacker_ram_3 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_54_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_kernel_unpacker_ram_3;
architecture structural of mh_72_bit_kernel_unpacker_ram_3 is 
  signal slice_71_down_to_54_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_35_down_to_18_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal data_delay_5_q_net : std_logic;
  signal slice_53_down_to_36_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal data_delay_4_q_net : std_logic;
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal slice_71_down_to_54_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_6_q_net : std_logic;
  signal data_delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_point_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_2_full_net : std_logic;
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_2_empty_net : std_logic;
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_2_op_net : std_logic_vector( 2-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal zero_out_op_net : std_logic_vector( 72-1 downto 0 );
  signal store_in_fifo_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 2-1 downto 0 );
begin
  x71_downto_54_fifo_0 <= slice_71_down_to_54_y_net;
  x53_downto_36_fifo_0 <= slice_53_down_to_36_y_net;
  x35_downto_18_fifo_0 <= slice_35_down_to_18_y_net;
  x17_downto_0_fifo_0 <= slice_17_down_to_0_y_net;
  x71_downto_54_fifo_1 <= slice_71_down_to_54_y_net_x0;
  x53_downto_36_fifo_1 <= slice_53_down_to_36_y_net_x0;
  x35_downto_18_fifo_1 <= slice_35_down_to_18_y_net_x0;
  x17_downto_0_fifo_1 <= slice_17_down_to_0_y_net_x0;
  x71_downto_54_fifo_2 <= slice_71_down_to_54_y_net_x1;
  x53_downto_36_fifo_2 <= slice_53_down_to_36_y_net_x1;
  x35_downto_18_fifo_2 <= slice_35_down_to_18_y_net_x1;
  x17_downto_0_fifo_2 <= slice_17_down_to_0_y_net_x1;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_3_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_kernel_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_0_x2 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net,
    x53_downto_36 => slice_53_down_to_36_y_net,
    x35_downto_18 => slice_35_down_to_18_y_net,
    x17_downto_0 => slice_17_down_to_0_y_net
  );
  unpack_kernel_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_1_x2 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x0,
    x53_downto_36 => slice_53_down_to_36_y_net_x0,
    x35_downto_18 => slice_35_down_to_18_y_net_x0,
    x17_downto_0 => slice_17_down_to_0_y_net_x0
  );
  unpack_kernel_72_bit_fifo_2 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_2_x2 
  port map (
    x72_bit_input => x72bit_frame_fifo_2_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x1,
    x53_downto_36 => slice_53_down_to_36_y_net_x1,
    x35_downto_18 => slice_35_down_to_18_y_net_x1,
    x17_downto_0 => slice_17_down_to_0_y_net_x1
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_delay_3_q_net,
    we => data_delay_4_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_5_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  x72bit_frame_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_6_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_2_dout_net,
    empty => x72bit_frame_fifo_2_empty_net,
    full => x72bit_frame_fifo_2_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_0_q_net
  );
  data_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_1_q_net
  );
  data_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_2_q_net
  );
  data_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_3_q_net
  );
  data_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_4_q_net
  );
  data_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_5_q_net
  );
  data_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_6_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  fifo_2 : entity xil_defaultlib.sysgen_constant_9d2d62a34e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_2_op_net
  );
  last_point_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => last_point_delay_q_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => last_point_delay_q_net,
    d1 => store_in_fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_bypass_fifo_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_2_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_2_y_net
  );
  logical : entity xil_defaultlib.sysgen_logical_17bd555d9a 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_1_empty_net,
    d1(0) => x72bit_frame_fifo_2_empty_net,
    d2(0) => x72bit_frame_fifo_0_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  store_in_fifo_2 : entity xil_defaultlib.sysgen_relational_bf21415019 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_2_op_net
  );
  sync_frame_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  write_to_fifo_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_2_y_net
  );
  zero_out : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_out_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => data_delay_2_q_net,
    d1 => zero_out_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 4/Unpack Kernel 72 Bit FIFO 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_0_x3 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_0_x3;
architecture structural of mh_unpack_kernel_72_bit_fifo_0_x3 is 
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_0_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_0_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 4/Unpack Kernel 72 Bit FIFO 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_1_x3 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_1_x3;
architecture structural of mh_unpack_kernel_72_bit_fifo_1_x3 is 
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_1_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_1_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 4/Unpack Kernel 72 Bit FIFO 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_unpack_kernel_72_bit_fifo_2_x3 is
  port (
    x72_bit_input : in std_logic_vector( 72-1 downto 0 );
    x71_downto_54 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_unpack_kernel_72_bit_fifo_2_x3;
architecture structural of mh_unpack_kernel_72_bit_fifo_2_x3 is 
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
begin
  x71_downto_54 <= slice_71_down_to_54_y_net;
  x53_downto_36 <= slice_53_down_to_36_y_net;
  x35_downto_18 <= slice_35_down_to_18_y_net;
  x17_downto_0 <= slice_17_down_to_0_y_net;
  x72bit_frame_fifo_2_dout_net <= x72_bit_input;
  slice_17_down_to_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_17_down_to_0_y_net
  );
  slice_35_down_to_18 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_35_down_to_18_y_net
  );
  slice_53_down_to_36 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 36,
    new_msb => 53,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_53_down_to_36_y_net
  );
  slice_71_down_to_54 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 54,
    new_msb => 71,
    x_width => 72,
    y_width => 18
  )
  port map (
    x => x72bit_frame_fifo_2_dout_net,
    y => slice_71_down_to_54_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/72 Bit Kernel Unpacker RAM 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_72_bit_kernel_unpacker_ram_4 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    enable : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    last_point : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x71_downto_54_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_0 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_1 : out std_logic_vector( 18-1 downto 0 );
    x71_downto_54_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x53_downto_36_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x35_downto_18_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    x17_downto_0_fifo_2 : out std_logic_vector( 18-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_a_fifo : out std_logic_vector( 1-1 downto 0 )
  );
end mh_72_bit_kernel_unpacker_ram_4;
architecture structural of mh_72_bit_kernel_unpacker_ram_4 is 
  signal store_in_fifo_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal sync_frame_counter_op_net : std_logic_vector( 2-1 downto 0 );
  signal last_value_bypass_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal zero_out_op_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_2_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_53_down_to_36_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal data_in_delay_1_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_0_dout_net : std_logic_vector( 72-1 downto 0 );
  signal slice_53_down_to_36_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x72bit_frame_fifo_1_dout_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_empty_net : std_logic;
  signal data_delay_4_q_net : std_logic;
  signal clk_net : std_logic;
  signal slice_17_down_to_0_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal data_delay_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal x72bit_frame_fifo_0_full_net : std_logic;
  signal slice_35_down_to_18_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal bypass_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_2_full_net : std_logic;
  signal data_delay_5_q_net : std_logic;
  signal x72bit_frame_fifo_1_empty_net : std_logic;
  signal enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_1_full_net : std_logic;
  signal bypass_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_6_q_net : std_logic;
  signal bypass_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal zero_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal data_delay_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_point_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal x72bit_frame_fifo_2_empty_net : std_logic;
  signal write_to_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal data_delay_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal fifo_2_op_net : std_logic_vector( 2-1 downto 0 );
  signal fifo_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_to_fifo_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal store_in_fifo_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_bypass_fifo_0_y_net : std_logic_vector( 1-1 downto 0 );
begin
  x71_downto_54_fifo_0 <= slice_71_down_to_54_y_net;
  x53_downto_36_fifo_0 <= slice_53_down_to_36_y_net;
  x35_downto_18_fifo_0 <= slice_35_down_to_18_y_net;
  x17_downto_0_fifo_0 <= slice_17_down_to_0_y_net;
  x71_downto_54_fifo_1 <= slice_71_down_to_54_y_net_x0;
  x53_downto_36_fifo_1 <= slice_53_down_to_36_y_net_x0;
  x35_downto_18_fifo_1 <= slice_35_down_to_18_y_net_x0;
  x17_downto_0_fifo_1 <= slice_17_down_to_0_y_net_x0;
  x71_downto_54_fifo_2 <= slice_71_down_to_54_y_net_x1;
  x53_downto_36_fifo_2 <= slice_53_down_to_36_y_net_x1;
  x35_downto_18_fifo_2 <= slice_35_down_to_18_y_net_x1;
  x17_downto_0_fifo_2 <= slice_17_down_to_0_y_net_x1;
  valid_out <= valid_q_net;
  wrote_to_a_fifo <= logical_y_net;
  data_in_delay_1_ram_4_q_net <= data_in;
  valid_delay_1_q_net <= enable;
  read_out_y_net <= read_enable;
  last_value_enable_y_net <= last_point;
  clk_net <= clk_1;
  ce_net <= ce_1;
  unpack_kernel_72_bit_fifo_0 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_0_x3 
  port map (
    x72_bit_input => x72bit_frame_fifo_0_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net,
    x53_downto_36 => slice_53_down_to_36_y_net,
    x35_downto_18 => slice_35_down_to_18_y_net,
    x17_downto_0 => slice_17_down_to_0_y_net
  );
  unpack_kernel_72_bit_fifo_1 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_1_x3 
  port map (
    x72_bit_input => x72bit_frame_fifo_1_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x0,
    x53_downto_36 => slice_53_down_to_36_y_net_x0,
    x35_downto_18 => slice_35_down_to_18_y_net_x0,
    x17_downto_0 => slice_17_down_to_0_y_net_x0
  );
  unpack_kernel_72_bit_fifo_2 : entity xil_defaultlib.mh_unpack_kernel_72_bit_fifo_2_x3 
  port map (
    x72_bit_input => x72bit_frame_fifo_2_dout_net,
    x71_downto_54 => slice_71_down_to_54_y_net_x1,
    x53_downto_36 => slice_53_down_to_36_y_net_x1,
    x35_downto_18 => slice_35_down_to_18_y_net_x1,
    x17_downto_0 => slice_17_down_to_0_y_net_x1
  );
  x72bit_frame_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => data_delay_3_q_net,
    we => data_delay_4_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_0_dout_net,
    empty => x72bit_frame_fifo_0_empty_net,
    full => x72bit_frame_fifo_0_full_net
  );
  x72bit_frame_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_5_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_1_dout_net,
    empty => x72bit_frame_fifo_1_empty_net,
    full => x72bit_frame_fifo_1_full_net
  );
  x72bit_frame_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i0",
    data_count_width => 4,
    data_width => 72,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => zero_value_y_net,
    we => data_delay_6_q_net,
    re => read_out_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => x72bit_frame_fifo_2_dout_net,
    empty => x72bit_frame_fifo_2_empty_net,
    full => x72bit_frame_fifo_2_full_net
  );
  bypass_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay_q_net
  );
  bypass_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay1_q_net
  );
  bypass_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => bypass_delay2_q_net
  );
  data_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_1_ram_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_0_q_net
  );
  data_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_1_q_net
  );
  data_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_2_q_net
  );
  data_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_delay_3_q_net
  );
  data_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_4_q_net
  );
  data_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_5_q_net
  );
  data_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_to_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q(0) => data_delay_6_q_net
  );
  enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay_q_net
  );
  fifo_0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_0_op_net
  );
  fifo_1 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_1_op_net
  );
  fifo_2 : entity xil_defaultlib.sysgen_constant_9d2d62a34e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => fifo_2_op_net
  );
  last_point_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_value_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    q => last_point_delay_q_net
  );
  last_value_bypass_fifo_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => last_point_delay_q_net,
    d1 => store_in_fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_0_y_net
  );
  last_value_bypass_fifo_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_1_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_1_y_net
  );
  last_value_bypass_fifo_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => store_in_fifo_2_op_net,
    d1 => last_point_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_bypass_fifo_2_y_net
  );
  logical : entity xil_defaultlib.sysgen_logical_17bd555d9a 
  port map (
    clr => '0',
    d0(0) => x72bit_frame_fifo_0_empty_net,
    d1(0) => x72bit_frame_fifo_1_empty_net,
    d2(0) => x72bit_frame_fifo_2_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  store_in_fifo_0 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_0_op_net
  );
  store_in_fifo_1 : entity xil_defaultlib.sysgen_relational_4dac6f3791 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_1_op_net
  );
  store_in_fifo_2 : entity xil_defaultlib.sysgen_relational_bf21415019 
  port map (
    clr => '0',
    a => sync_frame_counter_op_net,
    b => fifo_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => store_in_fifo_2_op_net
  );
  sync_frame_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => last_value_enable_y_net,
    en => valid_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => sync_frame_counter_op_net
  );
  valid : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => read_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_q_net
  );
  write_to_fifo_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => last_value_bypass_fifo_0_y_net,
    d1 => bypass_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_0_y_net
  );
  write_to_fifo_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_1_y_net
  );
  write_to_fifo_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => bypass_delay_q_net,
    d1 => last_value_bypass_fifo_2_y_net,
    clk => clk_net,
    ce => ce_net,
    y => write_to_fifo_2_y_net
  );
  zero_out : entity xil_defaultlib.sysgen_constant_fcb4de174e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_out_op_net
  );
  zero_value : entity xil_defaultlib.sysgen_mux_f33d45cf5b 
  port map (
    clr => '0',
    sel => bypass_delay2_q_net,
    d0 => data_delay_2_q_net,
    d1 => zero_out_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer/Data Point Tracker
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_data_point_tracker_x0 is
  port (
    data_in_ram_0 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_1 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_2 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_3 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_4 : in std_logic_vector( 72-1 downto 0 );
    valid_enable_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_out_ram_0 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_1 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_2 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_3 : out std_logic_vector( 72-1 downto 0 );
    data_out_ram_4 : out std_logic_vector( 72-1 downto 0 );
    valid_enable_out : out std_logic_vector( 1-1 downto 0 );
    last_value_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_data_point_tracker_x0;
architecture structural of mh_data_point_tracker_x0 is 
  signal data_in_delay_1_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_0_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
  signal clk_net : std_logic;
  signal data_in_delay_1_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal data_in_delay_0_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_1_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_point_counter_op_net : std_logic_vector( 7-1 downto 0 );
  signal data_in_delay_0_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_data_point_value_op_net : std_logic_vector( 7-1 downto 0 );
  signal data_in_delay_0_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal data_in_delay_0_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal last_point_op_net : std_logic_vector( 1-1 downto 0 );
  signal valid_delay_0_q_net : std_logic_vector( 1-1 downto 0 );
begin
  data_out_ram_0 <= data_in_delay_1_ram_0_q_net;
  data_out_ram_1 <= data_in_delay_1_ram_1_q_net;
  data_out_ram_2 <= data_in_delay_1_ram_2_q_net;
  data_out_ram_3 <= data_in_delay_1_ram_3_q_net;
  data_out_ram_4 <= data_in_delay_1_ram_4_q_net;
  valid_enable_out <= valid_delay_1_q_net;
  last_value_out <= last_value_enable_y_net;
  dual_port_ram_0_douta_net <= data_in_ram_0;
  dual_port_ram_1_douta_net <= data_in_ram_1;
  dual_port_ram_2_douta_net <= data_in_ram_2;
  dual_port_ram_3_douta_net <= data_in_ram_3;
  dual_port_ram_4_douta_net <= data_in_ram_4;
  convert_to_bool_dout_net <= valid_enable_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  data_in_delay_0_ram_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_0_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_0_q_net
  );
  data_in_delay_0_ram_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_1_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_1_q_net
  );
  data_in_delay_0_ram_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_2_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_2_q_net
  );
  data_in_delay_0_ram_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_3_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_3_q_net
  );
  data_in_delay_0_ram_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => dual_port_ram_4_douta_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_0_ram_4_q_net
  );
  data_in_delay_1_ram_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_0_q_net
  );
  data_in_delay_1_ram_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_1_q_net
  );
  data_in_delay_1_ram_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_2_q_net
  );
  data_in_delay_1_ram_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_3_q_net
  );
  data_in_delay_1_ram_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_delay_0_ram_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_in_delay_1_ram_4_q_net
  );
  data_point_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 99,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i0",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    rst => "0",
    clr => '0',
    en => convert_to_bool_dout_net,
    clk => clk_net,
    ce => ce_net,
    op => data_point_counter_op_net
  );
  last_data_point_value : entity xil_defaultlib.sysgen_constant_b4f986d24f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => last_data_point_value_op_net
  );
  last_point : entity xil_defaultlib.sysgen_relational_d18eb5aea1 
  port map (
    clr => '0',
    a => data_point_counter_op_net,
    b => last_data_point_value_op_net,
    clk => clk_net,
    ce => ce_net,
    op => last_point_op_net
  );
  last_value_enable : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => valid_delay_0_q_net,
    d1 => last_point_op_net,
    clk => clk_net,
    ce => ce_net,
    y => last_value_enable_y_net
  );
  valid_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_to_bool_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_delay_0_q_net
  );
  valid_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_delay_1_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Kernel RAM Slicer
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_ram_slicer is
  port (
    kernel_data_in_ram_0 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_1 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_2 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_3 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_4 : in std_logic_vector( 72-1 downto 0 );
    valid_in : in std_logic_vector( 1-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11_ram_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_0_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11_ram_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_0_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11_ram_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_0_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11_ram_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_0_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10_ram_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11_ram_4 : out std_logic_vector( 18-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_0 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_1 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_2 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_3 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_ram_4 : out std_logic_vector( 1-1 downto 0 );
    wrote_to_last_fifo_trigger : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_ram_slicer;
architecture structural of mh_kernel_ram_slicer is 
  signal delay_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal valid_sync_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_54_y_net_x13 : std_logic_vector( 18-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice_53_down_to_36_y_net_x13 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x13 : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal slice_53_down_to_36_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal slice_17_down_to_0_y_net_x13 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal last_fifo_written_to_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_54_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal data_in_delay_1_ram_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_18_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal data_in_delay_1_ram_2_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_18_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net : std_logic_vector( 18-1 downto 0 );
  signal last_value_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice_35_down_to_18_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice_17_down_to_0_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal valid_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal slice_53_down_to_36_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_71_down_to_54_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal data_in_delay_1_ram_1_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_71_down_to_54_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal data_in_delay_1_ram_3_q_net : std_logic_vector( 72-1 downto 0 );
  signal slice_35_down_to_18_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal valid_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice_53_down_to_36_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal slice_35_down_to_18_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_17_down_to_0_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal slice_71_down_to_54_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_53_down_to_36_y_net : std_logic_vector( 18-1 downto 0 );
  signal data_in_delay_1_ram_4_q_net : std_logic_vector( 72-1 downto 0 );
begin
  kernel_18_bit_value_0_ram_0 <= delay_3_q_net;
  kernel_18_bit_value_1_ram_0 <= delay_2_q_net;
  kernel_18_bit_value_2_ram_0 <= delay_1_q_net;
  kernel_18_bit_value_3_ram_0 <= delay_0_q_net;
  kernel_18_bit_value_4_ram_0 <= delay_7_q_net;
  kernel_18_bit_value_5_ram_0 <= delay_6_q_net;
  kernel_18_bit_value_6_ram_0 <= delay_5_q_net;
  kernel_18_bit_value_7_ram_0 <= delay_4_q_net;
  kernel_18_bit_value_8_ram_0 <= delay_11_q_net;
  kernel_18_bit_value_9_ram_0 <= delay_10_q_net;
  kernel_18_bit_value_10_ram_0 <= delay_9_q_net;
  kernel_18_bit_value_11_ram_0 <= delay_8_q_net;
  kernel_18_bit_value_0_ram_1 <= delay_17_q_net;
  kernel_18_bit_value_1_ram_1 <= delay_16_q_net;
  kernel_18_bit_value_2_ram_1 <= delay_13_q_net;
  kernel_18_bit_value_3_ram_1 <= delay_12_q_net;
  kernel_18_bit_value_4_ram_1 <= delay_21_q_net;
  kernel_18_bit_value_5_ram_1 <= delay_20_q_net;
  kernel_18_bit_value_6_ram_1 <= delay_19_q_net;
  kernel_18_bit_value_7_ram_1 <= delay_18_q_net;
  kernel_18_bit_value_8_ram_1 <= delay_15_q_net;
  kernel_18_bit_value_9_ram_1 <= delay_14_q_net;
  kernel_18_bit_value_10_ram_1 <= delay_23_q_net;
  kernel_18_bit_value_11_ram_1 <= delay_22_q_net;
  kernel_18_bit_value_0_ram_2 <= delay_29_q_net;
  kernel_18_bit_value_1_ram_2 <= delay_28_q_net;
  kernel_18_bit_value_2_ram_2 <= delay_25_q_net;
  kernel_18_bit_value_3_ram_2 <= delay_24_q_net;
  kernel_18_bit_value_4_ram_2 <= delay_33_q_net;
  kernel_18_bit_value_5_ram_2 <= delay_32_q_net;
  kernel_18_bit_value_6_ram_2 <= delay_31_q_net;
  kernel_18_bit_value_7_ram_2 <= delay_30_q_net;
  kernel_18_bit_value_8_ram_2 <= delay_27_q_net;
  kernel_18_bit_value_9_ram_2 <= delay_26_q_net;
  kernel_18_bit_value_10_ram_2 <= delay_35_q_net;
  kernel_18_bit_value_11_ram_2 <= delay_34_q_net;
  kernel_18_bit_value_0_ram_3 <= delay_41_q_net;
  kernel_18_bit_value_1_ram_3 <= delay_40_q_net;
  kernel_18_bit_value_2_ram_3 <= delay_37_q_net;
  kernel_18_bit_value_3_ram_3 <= delay_36_q_net;
  kernel_18_bit_value_4_ram_3 <= delay_45_q_net;
  kernel_18_bit_value_5_ram_3 <= delay_44_q_net;
  kernel_18_bit_value_6_ram_3 <= delay_43_q_net;
  kernel_18_bit_value_7_ram_3 <= delay_42_q_net;
  kernel_18_bit_value_8_ram_3 <= delay_39_q_net;
  kernel_18_bit_value_9_ram_3 <= delay_38_q_net;
  kernel_18_bit_value_10_ram_3 <= delay_47_q_net;
  kernel_18_bit_value_11_ram_3 <= delay_46_q_net;
  kernel_18_bit_value_0_ram_4 <= delay_53_q_net;
  kernel_18_bit_value_1_ram_4 <= delay_52_q_net;
  kernel_18_bit_value_2_ram_4 <= delay_49_q_net;
  kernel_18_bit_value_3_ram_4 <= delay_48_q_net;
  kernel_18_bit_value_4_ram_4 <= delay_57_q_net;
  kernel_18_bit_value_5_ram_4 <= delay_56_q_net;
  kernel_18_bit_value_6_ram_4 <= delay_55_q_net;
  kernel_18_bit_value_7_ram_4 <= delay_54_q_net;
  kernel_18_bit_value_8_ram_4 <= delay_51_q_net;
  kernel_18_bit_value_9_ram_4 <= delay_50_q_net;
  kernel_18_bit_value_10_ram_4 <= delay_59_q_net;
  kernel_18_bit_value_11_ram_4 <= delay_58_q_net;
  valid_out <= valid_sync_y_net;
  wrote_to_last_fifo_ram_0 <= logical_y_net_x3;
  wrote_to_last_fifo_ram_1 <= logical_y_net_x2;
  wrote_to_last_fifo_ram_2 <= logical_y_net_x1;
  wrote_to_last_fifo_ram_3 <= logical_y_net_x0;
  wrote_to_last_fifo_ram_4 <= logical_y_net;
  wrote_to_last_fifo_trigger <= last_fifo_written_to_1_q_net;
  dual_port_ram_0_douta_net <= kernel_data_in_ram_0;
  dual_port_ram_1_douta_net <= kernel_data_in_ram_1;
  dual_port_ram_2_douta_net <= kernel_data_in_ram_2;
  dual_port_ram_3_douta_net <= kernel_data_in_ram_3;
  dual_port_ram_4_douta_net <= kernel_data_in_ram_4;
  convert_to_bool_dout_net <= valid_in;
  read_out_y_net <= read_enable;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x72_bit_kernel_unpacker_ram_0 : entity xil_defaultlib.mh_72_bit_kernel_unpacker_ram_0 
  port map (
    data_in => data_in_delay_1_ram_0_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_54_fifo_0 => slice_71_down_to_54_y_net_x13,
    x53_downto_36_fifo_0 => slice_53_down_to_36_y_net_x13,
    x35_downto_18_fifo_0 => slice_35_down_to_18_y_net_x13,
    x17_downto_0_fifo_0 => slice_17_down_to_0_y_net_x13,
    x71_downto_54_fifo_1 => slice_71_down_to_54_y_net_x12,
    x53_downto_36_fifo_1 => slice_53_down_to_36_y_net_x12,
    x35_downto_18_fifo_1 => slice_35_down_to_18_y_net_x12,
    x17_downto_0_fifo_1 => slice_17_down_to_0_y_net_x12,
    x71_downto_54_fifo_2 => slice_71_down_to_54_y_net_x11,
    x53_downto_36_fifo_2 => slice_53_down_to_36_y_net_x11,
    x35_downto_18_fifo_2 => slice_35_down_to_18_y_net_x11,
    x17_downto_0_fifo_2 => slice_17_down_to_0_y_net_x11,
    valid_out => valid_q_net_x3,
    wrote_to_a_fifo => logical_y_net_x3,
    wrote_to_last_fifo => last_fifo_written_to_1_q_net
  );
  x72_bit_kernel_unpacker_ram_1 : entity xil_defaultlib.mh_72_bit_kernel_unpacker_ram_1 
  port map (
    data_in => data_in_delay_1_ram_1_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_54_fifo_0 => slice_71_down_to_54_y_net_x10,
    x53_downto_36_fifo_0 => slice_53_down_to_36_y_net_x10,
    x35_downto_18_fifo_0 => slice_35_down_to_18_y_net_x10,
    x17_downto_0_fifo_0 => slice_17_down_to_0_y_net_x10,
    x71_downto_54_fifo_1 => slice_71_down_to_54_y_net_x9,
    x53_downto_36_fifo_1 => slice_53_down_to_36_y_net_x9,
    x35_downto_18_fifo_1 => slice_35_down_to_18_y_net_x9,
    x17_downto_0_fifo_1 => slice_17_down_to_0_y_net_x9,
    x71_downto_54_fifo_2 => slice_71_down_to_54_y_net_x8,
    x53_downto_36_fifo_2 => slice_53_down_to_36_y_net_x8,
    x35_downto_18_fifo_2 => slice_35_down_to_18_y_net_x8,
    x17_downto_0_fifo_2 => slice_17_down_to_0_y_net_x8,
    valid_out => valid_q_net_x2,
    wrote_to_a_fifo => logical_y_net_x2
  );
  x72_bit_kernel_unpacker_ram_2 : entity xil_defaultlib.mh_72_bit_kernel_unpacker_ram_2 
  port map (
    data_in => data_in_delay_1_ram_2_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_54_fifo_0 => slice_71_down_to_54_y_net_x7,
    x53_downto_36_fifo_0 => slice_53_down_to_36_y_net_x7,
    x35_downto_18_fifo_0 => slice_35_down_to_18_y_net_x7,
    x17_downto_0_fifo_0 => slice_17_down_to_0_y_net_x7,
    x71_downto_54_fifo_1 => slice_71_down_to_54_y_net_x6,
    x53_downto_36_fifo_1 => slice_53_down_to_36_y_net_x6,
    x35_downto_18_fifo_1 => slice_35_down_to_18_y_net_x6,
    x17_downto_0_fifo_1 => slice_17_down_to_0_y_net_x6,
    x71_downto_54_fifo_2 => slice_71_down_to_54_y_net_x5,
    x53_downto_36_fifo_2 => slice_53_down_to_36_y_net_x5,
    x35_downto_18_fifo_2 => slice_35_down_to_18_y_net_x5,
    x17_downto_0_fifo_2 => slice_17_down_to_0_y_net_x5,
    valid_out => valid_q_net_x1,
    wrote_to_a_fifo => logical_y_net_x1
  );
  x72_bit_kernel_unpacker_ram_3 : entity xil_defaultlib.mh_72_bit_kernel_unpacker_ram_3 
  port map (
    data_in => data_in_delay_1_ram_3_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_54_fifo_0 => slice_71_down_to_54_y_net_x4,
    x53_downto_36_fifo_0 => slice_53_down_to_36_y_net_x4,
    x35_downto_18_fifo_0 => slice_35_down_to_18_y_net_x4,
    x17_downto_0_fifo_0 => slice_17_down_to_0_y_net_x4,
    x71_downto_54_fifo_1 => slice_71_down_to_54_y_net_x3,
    x53_downto_36_fifo_1 => slice_53_down_to_36_y_net_x3,
    x35_downto_18_fifo_1 => slice_35_down_to_18_y_net_x3,
    x17_downto_0_fifo_1 => slice_17_down_to_0_y_net_x3,
    x71_downto_54_fifo_2 => slice_71_down_to_54_y_net_x2,
    x53_downto_36_fifo_2 => slice_53_down_to_36_y_net_x2,
    x35_downto_18_fifo_2 => slice_35_down_to_18_y_net_x2,
    x17_downto_0_fifo_2 => slice_17_down_to_0_y_net_x2,
    valid_out => valid_q_net_x0,
    wrote_to_a_fifo => logical_y_net_x0
  );
  x72_bit_kernel_unpacker_ram_4 : entity xil_defaultlib.mh_72_bit_kernel_unpacker_ram_4 
  port map (
    data_in => data_in_delay_1_ram_4_q_net,
    enable => valid_delay_1_q_net,
    read_enable => read_out_y_net,
    last_point => last_value_enable_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x71_downto_54_fifo_0 => slice_71_down_to_54_y_net_x1,
    x53_downto_36_fifo_0 => slice_53_down_to_36_y_net_x1,
    x35_downto_18_fifo_0 => slice_35_down_to_18_y_net_x1,
    x17_downto_0_fifo_0 => slice_17_down_to_0_y_net_x1,
    x71_downto_54_fifo_1 => slice_71_down_to_54_y_net_x0,
    x53_downto_36_fifo_1 => slice_53_down_to_36_y_net_x0,
    x35_downto_18_fifo_1 => slice_35_down_to_18_y_net_x0,
    x17_downto_0_fifo_1 => slice_17_down_to_0_y_net_x0,
    x71_downto_54_fifo_2 => slice_71_down_to_54_y_net,
    x53_downto_36_fifo_2 => slice_53_down_to_36_y_net,
    x35_downto_18_fifo_2 => slice_35_down_to_18_y_net,
    x17_downto_0_fifo_2 => slice_17_down_to_0_y_net,
    valid_out => valid_q_net,
    wrote_to_a_fifo => logical_y_net
  );
  data_point_tracker : entity xil_defaultlib.mh_data_point_tracker_x0 
  port map (
    data_in_ram_0 => dual_port_ram_0_douta_net,
    data_in_ram_1 => dual_port_ram_1_douta_net,
    data_in_ram_2 => dual_port_ram_2_douta_net,
    data_in_ram_3 => dual_port_ram_3_douta_net,
    data_in_ram_4 => dual_port_ram_4_douta_net,
    valid_enable_in => convert_to_bool_dout_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    data_out_ram_0 => data_in_delay_1_ram_0_q_net,
    data_out_ram_1 => data_in_delay_1_ram_1_q_net,
    data_out_ram_2 => data_in_delay_1_ram_2_q_net,
    data_out_ram_3 => data_in_delay_1_ram_3_q_net,
    data_out_ram_4 => data_in_delay_1_ram_4_q_net,
    valid_enable_out => valid_delay_1_q_net,
    last_value_out => last_value_enable_y_net
  );
  delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x13,
    clk => clk_net,
    ce => ce_net,
    q => delay_0_q_net
  );
  delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x13,
    clk => clk_net,
    ce => ce_net,
    q => delay_1_q_net
  );
  delay_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x11,
    clk => clk_net,
    ce => ce_net,
    q => delay_10_q_net
  );
  delay_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x11,
    clk => clk_net,
    ce => ce_net,
    q => delay_11_q_net
  );
  delay_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x10,
    clk => clk_net,
    ce => ce_net,
    q => delay_12_q_net
  );
  delay_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x10,
    clk => clk_net,
    ce => ce_net,
    q => delay_13_q_net
  );
  delay_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_14_q_net
  );
  delay_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_15_q_net
  );
  delay_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x10,
    clk => clk_net,
    ce => ce_net,
    q => delay_16_q_net
  );
  delay_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x10,
    clk => clk_net,
    ce => ce_net,
    q => delay_17_q_net
  );
  delay_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x9,
    clk => clk_net,
    ce => ce_net,
    q => delay_18_q_net
  );
  delay_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x9,
    clk => clk_net,
    ce => ce_net,
    q => delay_19_q_net
  );
  delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x13,
    clk => clk_net,
    ce => ce_net,
    q => delay_2_q_net
  );
  delay_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x9,
    clk => clk_net,
    ce => ce_net,
    q => delay_20_q_net
  );
  delay_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x9,
    clk => clk_net,
    ce => ce_net,
    q => delay_21_q_net
  );
  delay_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_22_q_net
  );
  delay_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_23_q_net
  );
  delay_24 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_24_q_net
  );
  delay_25 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_25_q_net
  );
  delay_26 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_26_q_net
  );
  delay_27 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_27_q_net
  );
  delay_28 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_28_q_net
  );
  delay_29 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_29_q_net
  );
  delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x13,
    clk => clk_net,
    ce => ce_net,
    q => delay_3_q_net
  );
  delay_30 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_30_q_net
  );
  delay_31 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_31_q_net
  );
  delay_32 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_32_q_net
  );
  delay_33 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_33_q_net
  );
  delay_34 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_34_q_net
  );
  delay_35 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_35_q_net
  );
  delay_36 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_36_q_net
  );
  delay_37 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_37_q_net
  );
  delay_38 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_38_q_net
  );
  delay_39 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_39_q_net
  );
  delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay_4_q_net
  );
  delay_40 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_40_q_net
  );
  delay_41 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_41_q_net
  );
  delay_42 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_42_q_net
  );
  delay_43 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_43_q_net
  );
  delay_44 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_44_q_net
  );
  delay_45 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_45_q_net
  );
  delay_46 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_46_q_net
  );
  delay_47 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_47_q_net
  );
  delay_48 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_48_q_net
  );
  delay_49 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_49_q_net
  );
  delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay_5_q_net
  );
  delay_50 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_50_q_net
  );
  delay_51 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_51_q_net
  );
  delay_52 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_52_q_net
  );
  delay_53 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_53_q_net
  );
  delay_54 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_54_q_net
  );
  delay_55 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_55_q_net
  );
  delay_56 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_56_q_net
  );
  delay_57 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_57_q_net
  );
  delay_58 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_58_q_net
  );
  delay_59 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_59_q_net
  );
  delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_35_down_to_18_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay_6_q_net
  );
  delay_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_17_down_to_0_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay_7_q_net
  );
  delay_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_71_down_to_54_y_net_x11,
    clk => clk_net,
    ce => ce_net,
    q => delay_8_q_net
  );
  delay_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => slice_53_down_to_36_y_net_x11,
    clk => clk_net,
    ce => ce_net,
    q => delay_9_q_net
  );
  valid_sync : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => valid_q_net_x3,
    d1 => valid_q_net_x2,
    d2 => valid_q_net_x1,
    d3 => valid_q_net_x0,
    d4 => valid_q_net,
    clk => clk_net,
    ce => ce_net,
    y => valid_sync_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem1/Delay Kernel Values RAM 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_0 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 12-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_delay_kernel_values_ram_0;
architecture structural of mh_delay_kernel_values_ram_0 is 
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 12-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_5_q_net <= frame_12_bit_bin_value_0;
  delay_4_q_net <= frame_12_bit_bin_value_1;
  delay_3_q_net <= frame_12_bit_bin_value_2;
  delay_2_q_net <= frame_12_bit_bin_value_3;
  delay_1_q_net <= frame_12_bit_bin_value_4;
  delay_0_q_net <= frame_12_bit_bin_value_5;
  delay_11_q_net <= frame_12_bit_bin_value_6;
  delay_10_q_net <= frame_12_bit_bin_value_7;
  delay_9_q_net <= frame_12_bit_bin_value_8;
  delay_8_q_net <= frame_12_bit_bin_value_9;
  delay_7_q_net <= frame_12_bit_bin_value_10;
  delay_6_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem1/Delay Kernel Values RAM 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_1 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 12-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_delay_kernel_values_ram_1;
architecture structural of mh_delay_kernel_values_ram_1 is 
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 12-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_19_q_net <= frame_12_bit_bin_value_0;
  delay_18_q_net <= frame_12_bit_bin_value_1;
  delay_17_q_net <= frame_12_bit_bin_value_2;
  delay_16_q_net <= frame_12_bit_bin_value_3;
  delay_13_q_net <= frame_12_bit_bin_value_4;
  delay_12_q_net <= frame_12_bit_bin_value_5;
  delay_15_q_net <= frame_12_bit_bin_value_6;
  delay_14_q_net <= frame_12_bit_bin_value_7;
  delay_23_q_net <= frame_12_bit_bin_value_8;
  delay_22_q_net <= frame_12_bit_bin_value_9;
  delay_21_q_net <= frame_12_bit_bin_value_10;
  delay_20_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem1/Delay Kernel Values RAM 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_2 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 12-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_delay_kernel_values_ram_2;
architecture structural of mh_delay_kernel_values_ram_2 is 
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 12-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_43_q_net <= frame_12_bit_bin_value_0;
  delay_42_q_net <= frame_12_bit_bin_value_1;
  delay_41_q_net <= frame_12_bit_bin_value_2;
  delay_36_q_net <= frame_12_bit_bin_value_3;
  delay_25_q_net <= frame_12_bit_bin_value_4;
  delay_24_q_net <= frame_12_bit_bin_value_5;
  delay_27_q_net <= frame_12_bit_bin_value_6;
  delay_26_q_net <= frame_12_bit_bin_value_7;
  delay_47_q_net <= frame_12_bit_bin_value_8;
  delay_46_q_net <= frame_12_bit_bin_value_9;
  delay_45_q_net <= frame_12_bit_bin_value_10;
  delay_44_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_42_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_44_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_36_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_26_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_46_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem1/Delay Kernel Values RAM 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_3 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 12-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_delay_kernel_values_ram_3;
architecture structural of mh_delay_kernel_values_ram_3 is 
  signal delay_29_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 12-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_35_q_net <= frame_12_bit_bin_value_0;
  delay_34_q_net <= frame_12_bit_bin_value_1;
  delay_33_q_net <= frame_12_bit_bin_value_2;
  delay_32_q_net <= frame_12_bit_bin_value_3;
  delay_29_q_net <= frame_12_bit_bin_value_4;
  delay_28_q_net <= frame_12_bit_bin_value_5;
  delay_31_q_net <= frame_12_bit_bin_value_6;
  delay_30_q_net <= frame_12_bit_bin_value_7;
  delay_40_q_net <= frame_12_bit_bin_value_8;
  delay_39_q_net <= frame_12_bit_bin_value_9;
  delay_38_q_net <= frame_12_bit_bin_value_10;
  delay_37_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_34_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_37_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_32_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_28_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_30_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_39_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem1/Delay Kernel Values RAM 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_4 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 12-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 12-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_delay_kernel_values_ram_4;
architecture structural of mh_delay_kernel_values_ram_4 is 
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 12-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_67_q_net <= frame_12_bit_bin_value_0;
  delay_66_q_net <= frame_12_bit_bin_value_1;
  delay_65_q_net <= frame_12_bit_bin_value_2;
  delay_60_q_net <= frame_12_bit_bin_value_3;
  delay_49_q_net <= frame_12_bit_bin_value_4;
  delay_48_q_net <= frame_12_bit_bin_value_5;
  delay_51_q_net <= frame_12_bit_bin_value_6;
  delay_50_q_net <= frame_12_bit_bin_value_7;
  delay_71_q_net <= frame_12_bit_bin_value_8;
  delay_70_q_net <= frame_12_bit_bin_value_9;
  delay_69_q_net <= frame_12_bit_bin_value_10;
  delay_68_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_66_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_68_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_60_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_48_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_50_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_70_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_subsystem1 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_12 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_13 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_14 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_15 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_16 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_17 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_18 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_19 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_20 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_21 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_22 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_23 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_24 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_25 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_26 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_27 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_28 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_29 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_30 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_31 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_32 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_33 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_34 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_35 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_36 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_37 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_38 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_39 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_40 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_41 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_42 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_43 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_44 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_45 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_46 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_47 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_48 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_49 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_50 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_51 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_52 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_53 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_54 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_55 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_56 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_57 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_58 : in std_logic_vector( 12-1 downto 0 );
    frame_12_bit_bin_value_59 : in std_logic_vector( 12-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    frame_12_bit_value_0 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_1 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_2 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_3 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_4 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_5 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_6 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_7 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_8 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_9 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_10 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_11 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_12 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_13 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_14 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_15 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_16 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_17 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_18 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_19 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_20 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_21 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_22 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_23 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_24 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_25 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_26 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_27 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_28 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_29 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_30 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_31 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_32 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_33 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_34 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_35 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_36 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_37 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_38 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_39 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_40 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_41 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_42 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_43 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_44 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_45 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_46 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_47 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_48 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_49 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_50 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_51 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_52 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_53 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_54 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_55 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_56 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_57 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_58 : out std_logic_vector( 12-1 downto 0 );
    frame_12_bit_value_59 : out std_logic_vector( 12-1 downto 0 )
  );
end mh_subsystem1;
architecture structural of mh_subsystem1 is 
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_67_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x1 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x2 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x2 : std_logic_vector( 12-1 downto 0 );
begin
  frame_12_bit_value_0 <= x12_bit_bin_value_0_q_net_x3;
  frame_12_bit_value_1 <= x12_bit_bin_value_1_q_net_x3;
  frame_12_bit_value_2 <= x12_bit_bin_value_2_q_net_x3;
  frame_12_bit_value_3 <= x12_bit_bin_value_3_q_net_x3;
  frame_12_bit_value_4 <= x12_bit_bin_value_4_q_net_x3;
  frame_12_bit_value_5 <= x12_bit_bin_value_5_q_net_x3;
  frame_12_bit_value_6 <= x12_bit_bin_value_6_q_net_x3;
  frame_12_bit_value_7 <= x12_bit_bin_value_7_q_net_x2;
  frame_12_bit_value_8 <= x12_bit_bin_value_8_q_net_x2;
  frame_12_bit_value_9 <= x12_bit_bin_value_9_q_net_x2;
  frame_12_bit_value_10 <= x12_bit_bin_value_10_q_net_x3;
  frame_12_bit_value_11 <= x12_bit_bin_value_11_q_net_x3;
  frame_12_bit_value_12 <= x12_bit_bin_value_0_q_net_x2;
  frame_12_bit_value_13 <= x12_bit_bin_value_1_q_net_x2;
  frame_12_bit_value_14 <= x12_bit_bin_value_2_q_net_x2;
  frame_12_bit_value_15 <= x12_bit_bin_value_3_q_net_x2;
  frame_12_bit_value_16 <= x12_bit_bin_value_4_q_net_x2;
  frame_12_bit_value_17 <= x12_bit_bin_value_5_q_net_x2;
  frame_12_bit_value_18 <= x12_bit_bin_value_6_q_net_x2;
  frame_12_bit_value_19 <= x12_bit_bin_value_7_q_net_x1;
  frame_12_bit_value_20 <= x12_bit_bin_value_8_q_net_x1;
  frame_12_bit_value_21 <= x12_bit_bin_value_9_q_net_x1;
  frame_12_bit_value_22 <= x12_bit_bin_value_10_q_net_x2;
  frame_12_bit_value_23 <= x12_bit_bin_value_11_q_net_x2;
  frame_12_bit_value_24 <= x12_bit_bin_value_0_q_net_x1;
  frame_12_bit_value_25 <= x12_bit_bin_value_1_q_net_x1;
  frame_12_bit_value_26 <= x12_bit_bin_value_2_q_net_x1;
  frame_12_bit_value_27 <= x12_bit_bin_value_3_q_net_x1;
  frame_12_bit_value_28 <= x12_bit_bin_value_4_q_net_x1;
  frame_12_bit_value_29 <= x12_bit_bin_value_5_q_net_x1;
  frame_12_bit_value_30 <= x12_bit_bin_value_6_q_net_x1;
  frame_12_bit_value_31 <= x12_bit_bin_value_7_q_net_x0;
  frame_12_bit_value_32 <= x12_bit_bin_value_8_q_net_x0;
  frame_12_bit_value_33 <= x12_bit_bin_value_9_q_net_x0;
  frame_12_bit_value_34 <= x12_bit_bin_value_10_q_net_x1;
  frame_12_bit_value_35 <= x12_bit_bin_value_11_q_net_x1;
  frame_12_bit_value_36 <= x12_bit_bin_value_0_q_net_x0;
  frame_12_bit_value_37 <= x12_bit_bin_value_1_q_net_x0;
  frame_12_bit_value_38 <= x12_bit_bin_value_2_q_net_x0;
  frame_12_bit_value_39 <= x12_bit_bin_value_3_q_net_x0;
  frame_12_bit_value_40 <= x12_bit_bin_value_4_q_net_x0;
  frame_12_bit_value_41 <= x12_bit_bin_value_5_q_net_x0;
  frame_12_bit_value_42 <= x12_bit_bin_value_6_q_net_x0;
  frame_12_bit_value_43 <= x12_bit_bin_value_7_q_net;
  frame_12_bit_value_44 <= x12_bit_bin_value_8_q_net;
  frame_12_bit_value_45 <= x12_bit_bin_value_9_q_net;
  frame_12_bit_value_46 <= x12_bit_bin_value_10_q_net_x0;
  frame_12_bit_value_47 <= x12_bit_bin_value_11_q_net_x0;
  frame_12_bit_value_48 <= x12_bit_bin_value_0_q_net;
  frame_12_bit_value_49 <= x12_bit_bin_value_1_q_net;
  frame_12_bit_value_50 <= x12_bit_bin_value_2_q_net;
  frame_12_bit_value_51 <= x12_bit_bin_value_3_q_net;
  frame_12_bit_value_52 <= x12_bit_bin_value_4_q_net;
  frame_12_bit_value_53 <= x12_bit_bin_value_5_q_net;
  frame_12_bit_value_54 <= x12_bit_bin_value_6_q_net;
  frame_12_bit_value_55 <= x12_bit_bin_value_7_q_net_x3;
  frame_12_bit_value_56 <= x12_bit_bin_value_8_q_net_x3;
  frame_12_bit_value_57 <= x12_bit_bin_value_9_q_net_x3;
  frame_12_bit_value_58 <= x12_bit_bin_value_10_q_net;
  frame_12_bit_value_59 <= x12_bit_bin_value_11_q_net;
  delay_5_q_net <= frame_12_bit_bin_value_0;
  delay_4_q_net <= frame_12_bit_bin_value_1;
  delay_3_q_net <= frame_12_bit_bin_value_2;
  delay_2_q_net <= frame_12_bit_bin_value_3;
  delay_1_q_net <= frame_12_bit_bin_value_4;
  delay_0_q_net <= frame_12_bit_bin_value_5;
  delay_11_q_net <= frame_12_bit_bin_value_6;
  delay_10_q_net <= frame_12_bit_bin_value_7;
  delay_9_q_net <= frame_12_bit_bin_value_8;
  delay_8_q_net <= frame_12_bit_bin_value_9;
  delay_7_q_net <= frame_12_bit_bin_value_10;
  delay_6_q_net <= frame_12_bit_bin_value_11;
  delay_19_q_net <= frame_12_bit_bin_value_12;
  delay_18_q_net <= frame_12_bit_bin_value_13;
  delay_17_q_net <= frame_12_bit_bin_value_14;
  delay_16_q_net <= frame_12_bit_bin_value_15;
  delay_13_q_net <= frame_12_bit_bin_value_16;
  delay_12_q_net <= frame_12_bit_bin_value_17;
  delay_15_q_net <= frame_12_bit_bin_value_18;
  delay_14_q_net <= frame_12_bit_bin_value_19;
  delay_23_q_net <= frame_12_bit_bin_value_20;
  delay_22_q_net <= frame_12_bit_bin_value_21;
  delay_21_q_net <= frame_12_bit_bin_value_22;
  delay_20_q_net <= frame_12_bit_bin_value_23;
  delay_43_q_net <= frame_12_bit_bin_value_24;
  delay_42_q_net <= frame_12_bit_bin_value_25;
  delay_41_q_net <= frame_12_bit_bin_value_26;
  delay_36_q_net <= frame_12_bit_bin_value_27;
  delay_25_q_net <= frame_12_bit_bin_value_28;
  delay_24_q_net <= frame_12_bit_bin_value_29;
  delay_27_q_net <= frame_12_bit_bin_value_30;
  delay_26_q_net <= frame_12_bit_bin_value_31;
  delay_47_q_net <= frame_12_bit_bin_value_32;
  delay_46_q_net <= frame_12_bit_bin_value_33;
  delay_45_q_net <= frame_12_bit_bin_value_34;
  delay_44_q_net <= frame_12_bit_bin_value_35;
  delay_35_q_net <= frame_12_bit_bin_value_36;
  delay_34_q_net <= frame_12_bit_bin_value_37;
  delay_33_q_net <= frame_12_bit_bin_value_38;
  delay_32_q_net <= frame_12_bit_bin_value_39;
  delay_29_q_net <= frame_12_bit_bin_value_40;
  delay_28_q_net <= frame_12_bit_bin_value_41;
  delay_31_q_net <= frame_12_bit_bin_value_42;
  delay_30_q_net <= frame_12_bit_bin_value_43;
  delay_40_q_net <= frame_12_bit_bin_value_44;
  delay_39_q_net <= frame_12_bit_bin_value_45;
  delay_38_q_net <= frame_12_bit_bin_value_46;
  delay_37_q_net <= frame_12_bit_bin_value_47;
  delay_67_q_net <= frame_12_bit_bin_value_48;
  delay_66_q_net <= frame_12_bit_bin_value_49;
  delay_65_q_net <= frame_12_bit_bin_value_50;
  delay_60_q_net <= frame_12_bit_bin_value_51;
  delay_49_q_net <= frame_12_bit_bin_value_52;
  delay_48_q_net <= frame_12_bit_bin_value_53;
  delay_51_q_net <= frame_12_bit_bin_value_54;
  delay_50_q_net <= frame_12_bit_bin_value_55;
  delay_71_q_net <= frame_12_bit_bin_value_56;
  delay_70_q_net <= frame_12_bit_bin_value_57;
  delay_69_q_net <= frame_12_bit_bin_value_58;
  delay_68_q_net <= frame_12_bit_bin_value_59;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay_kernel_values_ram_0 : entity xil_defaultlib.mh_delay_kernel_values_ram_0 
  port map (
    frame_12_bit_bin_value_0 => delay_5_q_net,
    frame_12_bit_bin_value_1 => delay_4_q_net,
    frame_12_bit_bin_value_2 => delay_3_q_net,
    frame_12_bit_bin_value_3 => delay_2_q_net,
    frame_12_bit_bin_value_4 => delay_1_q_net,
    frame_12_bit_bin_value_5 => delay_0_q_net,
    frame_12_bit_bin_value_6 => delay_11_q_net,
    frame_12_bit_bin_value_7 => delay_10_q_net,
    frame_12_bit_bin_value_8 => delay_9_q_net,
    frame_12_bit_bin_value_9 => delay_8_q_net,
    frame_12_bit_bin_value_10 => delay_7_q_net,
    frame_12_bit_bin_value_11 => delay_6_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x3,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x3,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x3,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x3,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x3,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x3,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x3,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x2,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x2,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x2,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x3,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x3
  );
  delay_kernel_values_ram_1 : entity xil_defaultlib.mh_delay_kernel_values_ram_1 
  port map (
    frame_12_bit_bin_value_0 => delay_19_q_net,
    frame_12_bit_bin_value_1 => delay_18_q_net,
    frame_12_bit_bin_value_2 => delay_17_q_net,
    frame_12_bit_bin_value_3 => delay_16_q_net,
    frame_12_bit_bin_value_4 => delay_13_q_net,
    frame_12_bit_bin_value_5 => delay_12_q_net,
    frame_12_bit_bin_value_6 => delay_15_q_net,
    frame_12_bit_bin_value_7 => delay_14_q_net,
    frame_12_bit_bin_value_8 => delay_23_q_net,
    frame_12_bit_bin_value_9 => delay_22_q_net,
    frame_12_bit_bin_value_10 => delay_21_q_net,
    frame_12_bit_bin_value_11 => delay_20_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x2,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x2,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x2,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x2,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x2,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x2,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x2,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x1,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x1,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x1,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x2,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x2
  );
  delay_kernel_values_ram_2 : entity xil_defaultlib.mh_delay_kernel_values_ram_2 
  port map (
    frame_12_bit_bin_value_0 => delay_43_q_net,
    frame_12_bit_bin_value_1 => delay_42_q_net,
    frame_12_bit_bin_value_2 => delay_41_q_net,
    frame_12_bit_bin_value_3 => delay_36_q_net,
    frame_12_bit_bin_value_4 => delay_25_q_net,
    frame_12_bit_bin_value_5 => delay_24_q_net,
    frame_12_bit_bin_value_6 => delay_27_q_net,
    frame_12_bit_bin_value_7 => delay_26_q_net,
    frame_12_bit_bin_value_8 => delay_47_q_net,
    frame_12_bit_bin_value_9 => delay_46_q_net,
    frame_12_bit_bin_value_10 => delay_45_q_net,
    frame_12_bit_bin_value_11 => delay_44_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x1,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x1,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x1,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x1,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x1,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x1,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x1,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x0,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x0,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x0,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x1,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x1
  );
  delay_kernel_values_ram_3 : entity xil_defaultlib.mh_delay_kernel_values_ram_3 
  port map (
    frame_12_bit_bin_value_0 => delay_35_q_net,
    frame_12_bit_bin_value_1 => delay_34_q_net,
    frame_12_bit_bin_value_2 => delay_33_q_net,
    frame_12_bit_bin_value_3 => delay_32_q_net,
    frame_12_bit_bin_value_4 => delay_29_q_net,
    frame_12_bit_bin_value_5 => delay_28_q_net,
    frame_12_bit_bin_value_6 => delay_31_q_net,
    frame_12_bit_bin_value_7 => delay_30_q_net,
    frame_12_bit_bin_value_8 => delay_40_q_net,
    frame_12_bit_bin_value_9 => delay_39_q_net,
    frame_12_bit_bin_value_10 => delay_38_q_net,
    frame_12_bit_bin_value_11 => delay_37_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x0,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x0,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x0,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x0,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x0,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x0,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x0,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x0,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x0
  );
  delay_kernel_values_ram_4 : entity xil_defaultlib.mh_delay_kernel_values_ram_4 
  port map (
    frame_12_bit_bin_value_0 => delay_67_q_net,
    frame_12_bit_bin_value_1 => delay_66_q_net,
    frame_12_bit_bin_value_2 => delay_65_q_net,
    frame_12_bit_bin_value_3 => delay_60_q_net,
    frame_12_bit_bin_value_4 => delay_49_q_net,
    frame_12_bit_bin_value_5 => delay_48_q_net,
    frame_12_bit_bin_value_6 => delay_51_q_net,
    frame_12_bit_bin_value_7 => delay_50_q_net,
    frame_12_bit_bin_value_8 => delay_71_q_net,
    frame_12_bit_bin_value_9 => delay_70_q_net,
    frame_12_bit_bin_value_10 => delay_69_q_net,
    frame_12_bit_bin_value_11 => delay_68_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x3,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x3,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x3,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem2/Delay Kernel Values RAM 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_0_x0 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_delay_kernel_values_ram_0_x0;
architecture structural of mh_delay_kernel_values_ram_0_x0 is 
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal delay_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 18-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_3_q_net <= frame_12_bit_bin_value_0;
  delay_2_q_net <= frame_12_bit_bin_value_1;
  delay_1_q_net <= frame_12_bit_bin_value_2;
  delay_0_q_net <= frame_12_bit_bin_value_3;
  delay_7_q_net <= frame_12_bit_bin_value_4;
  delay_6_q_net <= frame_12_bit_bin_value_5;
  delay_5_q_net <= frame_12_bit_bin_value_6;
  delay_4_q_net <= frame_12_bit_bin_value_7;
  delay_11_q_net <= frame_12_bit_bin_value_8;
  delay_10_q_net <= frame_12_bit_bin_value_9;
  delay_9_q_net <= frame_12_bit_bin_value_10;
  delay_8_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem2/Delay Kernel Values RAM 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_1_x0 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_delay_kernel_values_ram_1_x0;
architecture structural of mh_delay_kernel_values_ram_1_x0 is 
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 18-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_17_q_net <= frame_12_bit_bin_value_0;
  delay_16_q_net <= frame_12_bit_bin_value_1;
  delay_13_q_net <= frame_12_bit_bin_value_2;
  delay_12_q_net <= frame_12_bit_bin_value_3;
  delay_21_q_net <= frame_12_bit_bin_value_4;
  delay_20_q_net <= frame_12_bit_bin_value_5;
  delay_19_q_net <= frame_12_bit_bin_value_6;
  delay_18_q_net <= frame_12_bit_bin_value_7;
  delay_15_q_net <= frame_12_bit_bin_value_8;
  delay_14_q_net <= frame_12_bit_bin_value_9;
  delay_23_q_net <= frame_12_bit_bin_value_10;
  delay_22_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem2/Delay Kernel Values RAM 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_2_x0 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_delay_kernel_values_ram_2_x0;
architecture structural of mh_delay_kernel_values_ram_2_x0 is 
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_32_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 18-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_29_q_net <= frame_12_bit_bin_value_0;
  delay_28_q_net <= frame_12_bit_bin_value_1;
  delay_25_q_net <= frame_12_bit_bin_value_2;
  delay_24_q_net <= frame_12_bit_bin_value_3;
  delay_33_q_net <= frame_12_bit_bin_value_4;
  delay_32_q_net <= frame_12_bit_bin_value_5;
  delay_31_q_net <= frame_12_bit_bin_value_6;
  delay_30_q_net <= frame_12_bit_bin_value_7;
  delay_27_q_net <= frame_12_bit_bin_value_8;
  delay_26_q_net <= frame_12_bit_bin_value_9;
  delay_35_q_net <= frame_12_bit_bin_value_10;
  delay_34_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_28_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_34_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_32_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_30_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_26_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem2/Delay Kernel Values RAM 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_3_x0 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_delay_kernel_values_ram_3_x0;
architecture structural of mh_delay_kernel_values_ram_3_x0 is 
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 18-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_41_q_net <= frame_12_bit_bin_value_0;
  delay_40_q_net <= frame_12_bit_bin_value_1;
  delay_37_q_net <= frame_12_bit_bin_value_2;
  delay_36_q_net <= frame_12_bit_bin_value_3;
  delay_45_q_net <= frame_12_bit_bin_value_4;
  delay_44_q_net <= frame_12_bit_bin_value_5;
  delay_43_q_net <= frame_12_bit_bin_value_6;
  delay_42_q_net <= frame_12_bit_bin_value_7;
  delay_39_q_net <= frame_12_bit_bin_value_8;
  delay_38_q_net <= frame_12_bit_bin_value_9;
  delay_47_q_net <= frame_12_bit_bin_value_10;
  delay_46_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_46_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_37_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_36_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_44_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_42_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_39_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem2/Delay Kernel Values RAM 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_delay_kernel_values_ram_4_x0 is
  port (
    frame_12_bit_bin_value_0 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_1 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_2 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_3 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_4 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_5 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_6 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_7 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_8 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_9 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_10 : in std_logic_vector( 18-1 downto 0 );
    frame_12_bit_bin_value_11 : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_delay_kernel_values_ram_4_x0;
architecture structural of mh_delay_kernel_values_ram_4_x0 is 
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal x12_bit_bin_value_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_18_q_net : std_logic_vector( 18-1 downto 0 );
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net;
  delay_53_q_net <= frame_12_bit_bin_value_0;
  delay_52_q_net <= frame_12_bit_bin_value_1;
  delay_49_q_net <= frame_12_bit_bin_value_2;
  delay_48_q_net <= frame_12_bit_bin_value_3;
  delay_57_q_net <= frame_12_bit_bin_value_4;
  delay_56_q_net <= frame_12_bit_bin_value_5;
  delay_55_q_net <= frame_12_bit_bin_value_6;
  delay_54_q_net <= frame_12_bit_bin_value_7;
  delay_51_q_net <= frame_12_bit_bin_value_8;
  delay_50_q_net <= frame_12_bit_bin_value_9;
  delay_59_q_net <= frame_12_bit_bin_value_10;
  delay_58_q_net <= frame_12_bit_bin_value_11;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x12_bit_bin_value_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_0_q_net
  );
  x12_bit_bin_value_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_1_q_net
  );
  x12_bit_bin_value_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_10_q_net
  );
  x12_bit_bin_value_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_11_q_net
  );
  x12_bit_bin_value_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_12_q_net
  );
  x12_bit_bin_value_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_52_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_13_q_net
  );
  x12_bit_bin_value_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_14_q_net
  );
  x12_bit_bin_value_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_58_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_15_q_net
  );
  x12_bit_bin_value_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_16_q_net
  );
  x12_bit_bin_value_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_48_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_17_q_net
  );
  x12_bit_bin_value_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_18_q_net
  );
  x12_bit_bin_value_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_56_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_19_q_net
  );
  x12_bit_bin_value_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_2_q_net
  );
  x12_bit_bin_value_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_20_q_net
  );
  x12_bit_bin_value_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_54_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_21_q_net
  );
  x12_bit_bin_value_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_22_q_net
  );
  x12_bit_bin_value_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_50_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_23_q_net
  );
  x12_bit_bin_value_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_3_q_net
  );
  x12_bit_bin_value_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_4_q_net
  );
  x12_bit_bin_value_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_5_q_net
  );
  x12_bit_bin_value_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_6_q_net
  );
  x12_bit_bin_value_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_21_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_7_q_net
  );
  x12_bit_bin_value_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_8_q_net
  );
  x12_bit_bin_value_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_23_q_net,
    clk => clk_net,
    ce => ce_net,
    q => x12_bit_bin_value_9_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer/Subsystem2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_subsystem2 is
  port (
    kernel_18_bit_bin_value_0 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_1 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_2 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_3 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_4 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_5 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_6 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_7 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_8 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_9 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_10 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_11 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_12 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_13 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_14 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_15 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_16 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_17 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_18 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_19 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_20 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_21 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_22 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_23 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_24 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_25 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_26 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_27 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_28 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_29 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_30 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_31 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_32 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_33 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_34 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_35 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_36 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_37 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_38 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_39 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_40 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_41 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_42 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_43 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_44 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_45 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_46 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_47 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_48 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_49 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_50 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_51 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_52 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_53 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_54 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_55 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_56 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_57 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_58 : in std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_bin_value_59 : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_18_bit_value_0 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_2 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_3 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_4 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_5 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_6 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_7 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_8 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_9 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_10 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_11 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_12 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_13 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_14 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_15 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_16 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_17 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_18 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_19 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_20 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_21 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_22 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_23 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_24 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_25 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_26 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_27 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_28 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_29 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_30 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_31 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_32 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_33 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_34 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_35 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_36 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_37 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_38 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_39 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_40 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_41 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_42 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_43 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_44 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_45 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_46 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_47 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_48 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_49 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_50 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_51 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_52 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_53 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_54 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_55 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_56 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_57 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_58 : out std_logic_vector( 18-1 downto 0 );
    kernel_18_bit_value_59 : out std_logic_vector( 18-1 downto 0 )
  );
end mh_subsystem2;
architecture structural of mh_subsystem2 is 
  signal x12_bit_bin_value_1_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_58_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
begin
  kernel_18_bit_value_0 <= x12_bit_bin_value_0_q_net_x3;
  kernel_18_bit_value_1 <= x12_bit_bin_value_1_q_net_x3;
  kernel_18_bit_value_2 <= x12_bit_bin_value_2_q_net_x3;
  kernel_18_bit_value_3 <= x12_bit_bin_value_3_q_net_x3;
  kernel_18_bit_value_4 <= x12_bit_bin_value_4_q_net_x3;
  kernel_18_bit_value_5 <= x12_bit_bin_value_5_q_net_x3;
  kernel_18_bit_value_6 <= x12_bit_bin_value_6_q_net_x3;
  kernel_18_bit_value_7 <= x12_bit_bin_value_7_q_net_x2;
  kernel_18_bit_value_8 <= x12_bit_bin_value_8_q_net_x2;
  kernel_18_bit_value_9 <= x12_bit_bin_value_9_q_net_x2;
  kernel_18_bit_value_10 <= x12_bit_bin_value_10_q_net_x3;
  kernel_18_bit_value_11 <= x12_bit_bin_value_11_q_net_x3;
  kernel_18_bit_value_12 <= x12_bit_bin_value_0_q_net_x2;
  kernel_18_bit_value_13 <= x12_bit_bin_value_1_q_net_x2;
  kernel_18_bit_value_14 <= x12_bit_bin_value_2_q_net_x2;
  kernel_18_bit_value_15 <= x12_bit_bin_value_3_q_net_x2;
  kernel_18_bit_value_16 <= x12_bit_bin_value_4_q_net_x2;
  kernel_18_bit_value_17 <= x12_bit_bin_value_5_q_net_x2;
  kernel_18_bit_value_18 <= x12_bit_bin_value_6_q_net_x2;
  kernel_18_bit_value_19 <= x12_bit_bin_value_7_q_net_x1;
  kernel_18_bit_value_20 <= x12_bit_bin_value_8_q_net_x1;
  kernel_18_bit_value_21 <= x12_bit_bin_value_9_q_net_x1;
  kernel_18_bit_value_22 <= x12_bit_bin_value_10_q_net_x2;
  kernel_18_bit_value_23 <= x12_bit_bin_value_11_q_net_x2;
  kernel_18_bit_value_24 <= x12_bit_bin_value_0_q_net_x1;
  kernel_18_bit_value_25 <= x12_bit_bin_value_1_q_net_x1;
  kernel_18_bit_value_26 <= x12_bit_bin_value_2_q_net_x1;
  kernel_18_bit_value_27 <= x12_bit_bin_value_3_q_net_x1;
  kernel_18_bit_value_28 <= x12_bit_bin_value_4_q_net_x1;
  kernel_18_bit_value_29 <= x12_bit_bin_value_5_q_net_x1;
  kernel_18_bit_value_30 <= x12_bit_bin_value_6_q_net_x1;
  kernel_18_bit_value_31 <= x12_bit_bin_value_7_q_net_x0;
  kernel_18_bit_value_32 <= x12_bit_bin_value_8_q_net_x0;
  kernel_18_bit_value_33 <= x12_bit_bin_value_9_q_net_x0;
  kernel_18_bit_value_34 <= x12_bit_bin_value_10_q_net_x1;
  kernel_18_bit_value_35 <= x12_bit_bin_value_11_q_net_x1;
  kernel_18_bit_value_36 <= x12_bit_bin_value_0_q_net_x0;
  kernel_18_bit_value_37 <= x12_bit_bin_value_1_q_net_x0;
  kernel_18_bit_value_38 <= x12_bit_bin_value_2_q_net_x0;
  kernel_18_bit_value_39 <= x12_bit_bin_value_3_q_net_x0;
  kernel_18_bit_value_40 <= x12_bit_bin_value_4_q_net_x0;
  kernel_18_bit_value_41 <= x12_bit_bin_value_5_q_net_x0;
  kernel_18_bit_value_42 <= x12_bit_bin_value_6_q_net_x0;
  kernel_18_bit_value_43 <= x12_bit_bin_value_7_q_net;
  kernel_18_bit_value_44 <= x12_bit_bin_value_8_q_net;
  kernel_18_bit_value_45 <= x12_bit_bin_value_9_q_net;
  kernel_18_bit_value_46 <= x12_bit_bin_value_10_q_net_x0;
  kernel_18_bit_value_47 <= x12_bit_bin_value_11_q_net_x0;
  kernel_18_bit_value_48 <= x12_bit_bin_value_0_q_net;
  kernel_18_bit_value_49 <= x12_bit_bin_value_1_q_net;
  kernel_18_bit_value_50 <= x12_bit_bin_value_2_q_net;
  kernel_18_bit_value_51 <= x12_bit_bin_value_3_q_net;
  kernel_18_bit_value_52 <= x12_bit_bin_value_4_q_net;
  kernel_18_bit_value_53 <= x12_bit_bin_value_5_q_net;
  kernel_18_bit_value_54 <= x12_bit_bin_value_6_q_net;
  kernel_18_bit_value_55 <= x12_bit_bin_value_7_q_net_x3;
  kernel_18_bit_value_56 <= x12_bit_bin_value_8_q_net_x3;
  kernel_18_bit_value_57 <= x12_bit_bin_value_9_q_net_x3;
  kernel_18_bit_value_58 <= x12_bit_bin_value_10_q_net;
  kernel_18_bit_value_59 <= x12_bit_bin_value_11_q_net;
  delay_3_q_net <= kernel_18_bit_bin_value_0;
  delay_2_q_net <= kernel_18_bit_bin_value_1;
  delay_1_q_net <= kernel_18_bit_bin_value_2;
  delay_0_q_net <= kernel_18_bit_bin_value_3;
  delay_7_q_net <= kernel_18_bit_bin_value_4;
  delay_6_q_net <= kernel_18_bit_bin_value_5;
  delay_5_q_net <= kernel_18_bit_bin_value_6;
  delay_4_q_net <= kernel_18_bit_bin_value_7;
  delay_11_q_net <= kernel_18_bit_bin_value_8;
  delay_10_q_net <= kernel_18_bit_bin_value_9;
  delay_9_q_net <= kernel_18_bit_bin_value_10;
  delay_8_q_net <= kernel_18_bit_bin_value_11;
  delay_17_q_net <= kernel_18_bit_bin_value_12;
  delay_16_q_net <= kernel_18_bit_bin_value_13;
  delay_13_q_net <= kernel_18_bit_bin_value_14;
  delay_12_q_net <= kernel_18_bit_bin_value_15;
  delay_21_q_net <= kernel_18_bit_bin_value_16;
  delay_20_q_net <= kernel_18_bit_bin_value_17;
  delay_19_q_net <= kernel_18_bit_bin_value_18;
  delay_18_q_net <= kernel_18_bit_bin_value_19;
  delay_15_q_net <= kernel_18_bit_bin_value_20;
  delay_14_q_net <= kernel_18_bit_bin_value_21;
  delay_23_q_net <= kernel_18_bit_bin_value_22;
  delay_22_q_net <= kernel_18_bit_bin_value_23;
  delay_29_q_net <= kernel_18_bit_bin_value_24;
  delay_28_q_net <= kernel_18_bit_bin_value_25;
  delay_25_q_net <= kernel_18_bit_bin_value_26;
  delay_24_q_net <= kernel_18_bit_bin_value_27;
  delay_33_q_net <= kernel_18_bit_bin_value_28;
  delay_32_q_net <= kernel_18_bit_bin_value_29;
  delay_31_q_net <= kernel_18_bit_bin_value_30;
  delay_30_q_net <= kernel_18_bit_bin_value_31;
  delay_27_q_net <= kernel_18_bit_bin_value_32;
  delay_26_q_net <= kernel_18_bit_bin_value_33;
  delay_35_q_net <= kernel_18_bit_bin_value_34;
  delay_34_q_net <= kernel_18_bit_bin_value_35;
  delay_41_q_net <= kernel_18_bit_bin_value_36;
  delay_40_q_net <= kernel_18_bit_bin_value_37;
  delay_37_q_net <= kernel_18_bit_bin_value_38;
  delay_36_q_net <= kernel_18_bit_bin_value_39;
  delay_45_q_net <= kernel_18_bit_bin_value_40;
  delay_44_q_net <= kernel_18_bit_bin_value_41;
  delay_43_q_net <= kernel_18_bit_bin_value_42;
  delay_42_q_net <= kernel_18_bit_bin_value_43;
  delay_39_q_net <= kernel_18_bit_bin_value_44;
  delay_38_q_net <= kernel_18_bit_bin_value_45;
  delay_47_q_net <= kernel_18_bit_bin_value_46;
  delay_46_q_net <= kernel_18_bit_bin_value_47;
  delay_53_q_net <= kernel_18_bit_bin_value_48;
  delay_52_q_net <= kernel_18_bit_bin_value_49;
  delay_49_q_net <= kernel_18_bit_bin_value_50;
  delay_48_q_net <= kernel_18_bit_bin_value_51;
  delay_57_q_net <= kernel_18_bit_bin_value_52;
  delay_56_q_net <= kernel_18_bit_bin_value_53;
  delay_55_q_net <= kernel_18_bit_bin_value_54;
  delay_54_q_net <= kernel_18_bit_bin_value_55;
  delay_51_q_net <= kernel_18_bit_bin_value_56;
  delay_50_q_net <= kernel_18_bit_bin_value_57;
  delay_59_q_net <= kernel_18_bit_bin_value_58;
  delay_58_q_net <= kernel_18_bit_bin_value_59;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay_kernel_values_ram_0 : entity xil_defaultlib.mh_delay_kernel_values_ram_0_x0 
  port map (
    frame_12_bit_bin_value_0 => delay_3_q_net,
    frame_12_bit_bin_value_1 => delay_2_q_net,
    frame_12_bit_bin_value_2 => delay_1_q_net,
    frame_12_bit_bin_value_3 => delay_0_q_net,
    frame_12_bit_bin_value_4 => delay_7_q_net,
    frame_12_bit_bin_value_5 => delay_6_q_net,
    frame_12_bit_bin_value_6 => delay_5_q_net,
    frame_12_bit_bin_value_7 => delay_4_q_net,
    frame_12_bit_bin_value_8 => delay_11_q_net,
    frame_12_bit_bin_value_9 => delay_10_q_net,
    frame_12_bit_bin_value_10 => delay_9_q_net,
    frame_12_bit_bin_value_11 => delay_8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x3,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x3,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x3,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x3,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x3,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x3,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x3,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x2,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x2,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x2,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x3,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x3
  );
  delay_kernel_values_ram_1 : entity xil_defaultlib.mh_delay_kernel_values_ram_1_x0 
  port map (
    frame_12_bit_bin_value_0 => delay_17_q_net,
    frame_12_bit_bin_value_1 => delay_16_q_net,
    frame_12_bit_bin_value_2 => delay_13_q_net,
    frame_12_bit_bin_value_3 => delay_12_q_net,
    frame_12_bit_bin_value_4 => delay_21_q_net,
    frame_12_bit_bin_value_5 => delay_20_q_net,
    frame_12_bit_bin_value_6 => delay_19_q_net,
    frame_12_bit_bin_value_7 => delay_18_q_net,
    frame_12_bit_bin_value_8 => delay_15_q_net,
    frame_12_bit_bin_value_9 => delay_14_q_net,
    frame_12_bit_bin_value_10 => delay_23_q_net,
    frame_12_bit_bin_value_11 => delay_22_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x2,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x2,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x2,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x2,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x2,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x2,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x2,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x1,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x1,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x1,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x2,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x2
  );
  delay_kernel_values_ram_2 : entity xil_defaultlib.mh_delay_kernel_values_ram_2_x0 
  port map (
    frame_12_bit_bin_value_0 => delay_29_q_net,
    frame_12_bit_bin_value_1 => delay_28_q_net,
    frame_12_bit_bin_value_2 => delay_25_q_net,
    frame_12_bit_bin_value_3 => delay_24_q_net,
    frame_12_bit_bin_value_4 => delay_33_q_net,
    frame_12_bit_bin_value_5 => delay_32_q_net,
    frame_12_bit_bin_value_6 => delay_31_q_net,
    frame_12_bit_bin_value_7 => delay_30_q_net,
    frame_12_bit_bin_value_8 => delay_27_q_net,
    frame_12_bit_bin_value_9 => delay_26_q_net,
    frame_12_bit_bin_value_10 => delay_35_q_net,
    frame_12_bit_bin_value_11 => delay_34_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x1,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x1,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x1,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x1,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x1,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x1,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x1,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x0,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x0,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x0,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x1,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x1
  );
  delay_kernel_values_ram_3 : entity xil_defaultlib.mh_delay_kernel_values_ram_3_x0 
  port map (
    frame_12_bit_bin_value_0 => delay_41_q_net,
    frame_12_bit_bin_value_1 => delay_40_q_net,
    frame_12_bit_bin_value_2 => delay_37_q_net,
    frame_12_bit_bin_value_3 => delay_36_q_net,
    frame_12_bit_bin_value_4 => delay_45_q_net,
    frame_12_bit_bin_value_5 => delay_44_q_net,
    frame_12_bit_bin_value_6 => delay_43_q_net,
    frame_12_bit_bin_value_7 => delay_42_q_net,
    frame_12_bit_bin_value_8 => delay_39_q_net,
    frame_12_bit_bin_value_9 => delay_38_q_net,
    frame_12_bit_bin_value_10 => delay_47_q_net,
    frame_12_bit_bin_value_11 => delay_46_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x0,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x0,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x0,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x0,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x0,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x0,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x0,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x0,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x0
  );
  delay_kernel_values_ram_4 : entity xil_defaultlib.mh_delay_kernel_values_ram_4_x0 
  port map (
    frame_12_bit_bin_value_0 => delay_53_q_net,
    frame_12_bit_bin_value_1 => delay_52_q_net,
    frame_12_bit_bin_value_2 => delay_49_q_net,
    frame_12_bit_bin_value_3 => delay_48_q_net,
    frame_12_bit_bin_value_4 => delay_57_q_net,
    frame_12_bit_bin_value_5 => delay_56_q_net,
    frame_12_bit_bin_value_6 => delay_55_q_net,
    frame_12_bit_bin_value_7 => delay_54_q_net,
    frame_12_bit_bin_value_8 => delay_51_q_net,
    frame_12_bit_bin_value_9 => delay_50_q_net,
    frame_12_bit_bin_value_10 => delay_59_q_net,
    frame_12_bit_bin_value_11 => delay_58_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x3,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x3,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x3,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Data Slicer
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_data_slicer is
  port (
    data_in_ram_0 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_1 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_2 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_3 : in std_logic_vector( 72-1 downto 0 );
    data_in_ram_4 : in std_logic_vector( 72-1 downto 0 );
    frame_valid_in : in std_logic_vector( 1-1 downto 0 );
    kernel_data_in_ram_0 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_1 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_2 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_3 : in std_logic_vector( 72-1 downto 0 );
    kernel_data_in_ram_4 : in std_logic_vector( 72-1 downto 0 );
    kernel_valid_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    frame_pixel_0_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_1_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_2_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_3_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_4_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_5_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_6_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_7_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_8_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_9_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_10_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_11_at_offset_0 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_0_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_1_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_2_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_3_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_4_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_5_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_6_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_7_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_8_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_9_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_10_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_11_at_offset_1 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_0_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_1_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_2_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_3_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_4_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_5_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_6_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_7_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_8_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_9_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_10_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_11_at_offset_2 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_0_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_1_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_2_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_3_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_4_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_5_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_6_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_7_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_8_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_9_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_10_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_11_at_offset_3 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_0_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_1_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_2_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_3_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_4_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_5_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_6_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_7_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_8_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_9_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_10_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    frame_pixel_11_at_offset_4 : out std_logic_vector( 12-1 downto 0 );
    weight_0_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_1_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_2_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_3_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_4_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_5_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_6_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_7_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_8_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_9_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_10_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_11_at_offset_0 : out std_logic_vector( 18-1 downto 0 );
    weight_0_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_1_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_2_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_3_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_4_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_5_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_6_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_7_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_8_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_9_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_10_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_11_at_offset_1 : out std_logic_vector( 18-1 downto 0 );
    weight_0_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_1_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_2_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_3_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_4_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_5_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_6_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_7_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_8_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_9_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_10_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_11_at_offset_2 : out std_logic_vector( 18-1 downto 0 );
    weight_0_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_1_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_2_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_3_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_4_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_5_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_6_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_7_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_8_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_9_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_10_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_11_at_offset_3 : out std_logic_vector( 18-1 downto 0 );
    weight_0_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_1_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_2_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_3_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_4_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_5_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_6_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_7_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_8_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_9_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_10_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    weight_11_at_offset_4 : out std_logic_vector( 18-1 downto 0 );
    valid_data : out std_logic_vector( 1-1 downto 0 )
  );
end mh_data_slicer;
architecture structural of mh_data_slicer is 
  signal delay_51_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal valid_sync_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_44_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal read_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_33_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal logical_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 18-1 downto 0 );
  signal valid_sync_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_fifo_written_to_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 18-1 downto 0 );
  signal valid_out_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal data_valid_out_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_3_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal delay_4_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_4_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal convert_to_bool_dout_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_5_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal dual_port_ram_0_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_11_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal dual_port_ram_1_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal delay_3_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net_x0 : std_logic_vector( 12-1 downto 0 );
begin
  frame_pixel_0_at_offset_0 <= x12_bit_bin_value_0_q_net_x8;
  frame_pixel_1_at_offset_0 <= x12_bit_bin_value_1_q_net_x8;
  frame_pixel_2_at_offset_0 <= x12_bit_bin_value_2_q_net_x8;
  frame_pixel_3_at_offset_0 <= x12_bit_bin_value_3_q_net_x8;
  frame_pixel_4_at_offset_0 <= x12_bit_bin_value_4_q_net_x8;
  frame_pixel_5_at_offset_0 <= x12_bit_bin_value_5_q_net_x8;
  frame_pixel_6_at_offset_0 <= x12_bit_bin_value_6_q_net_x8;
  frame_pixel_7_at_offset_0 <= x12_bit_bin_value_7_q_net_x8;
  frame_pixel_8_at_offset_0 <= x12_bit_bin_value_8_q_net_x8;
  frame_pixel_9_at_offset_0 <= x12_bit_bin_value_9_q_net_x8;
  frame_pixel_10_at_offset_0 <= x12_bit_bin_value_10_q_net_x8;
  frame_pixel_11_at_offset_0 <= x12_bit_bin_value_11_q_net_x8;
  frame_pixel_0_at_offset_1 <= x12_bit_bin_value_0_q_net_x7;
  frame_pixel_1_at_offset_1 <= x12_bit_bin_value_1_q_net_x7;
  frame_pixel_2_at_offset_1 <= x12_bit_bin_value_2_q_net_x7;
  frame_pixel_3_at_offset_1 <= x12_bit_bin_value_3_q_net_x7;
  frame_pixel_4_at_offset_1 <= x12_bit_bin_value_4_q_net_x7;
  frame_pixel_5_at_offset_1 <= x12_bit_bin_value_5_q_net_x7;
  frame_pixel_6_at_offset_1 <= x12_bit_bin_value_6_q_net_x7;
  frame_pixel_7_at_offset_1 <= x12_bit_bin_value_7_q_net_x7;
  frame_pixel_8_at_offset_1 <= x12_bit_bin_value_8_q_net_x7;
  frame_pixel_9_at_offset_1 <= x12_bit_bin_value_9_q_net_x7;
  frame_pixel_10_at_offset_1 <= x12_bit_bin_value_10_q_net_x7;
  frame_pixel_11_at_offset_1 <= x12_bit_bin_value_11_q_net_x7;
  frame_pixel_0_at_offset_2 <= x12_bit_bin_value_0_q_net_x6;
  frame_pixel_1_at_offset_2 <= x12_bit_bin_value_1_q_net_x6;
  frame_pixel_2_at_offset_2 <= x12_bit_bin_value_2_q_net_x6;
  frame_pixel_3_at_offset_2 <= x12_bit_bin_value_3_q_net_x6;
  frame_pixel_4_at_offset_2 <= x12_bit_bin_value_4_q_net_x6;
  frame_pixel_5_at_offset_2 <= x12_bit_bin_value_5_q_net_x6;
  frame_pixel_6_at_offset_2 <= x12_bit_bin_value_6_q_net_x6;
  frame_pixel_7_at_offset_2 <= x12_bit_bin_value_7_q_net_x6;
  frame_pixel_8_at_offset_2 <= x12_bit_bin_value_8_q_net_x6;
  frame_pixel_9_at_offset_2 <= x12_bit_bin_value_9_q_net_x6;
  frame_pixel_10_at_offset_2 <= x12_bit_bin_value_10_q_net_x6;
  frame_pixel_11_at_offset_2 <= x12_bit_bin_value_11_q_net_x6;
  frame_pixel_0_at_offset_3 <= x12_bit_bin_value_0_q_net_x5;
  frame_pixel_1_at_offset_3 <= x12_bit_bin_value_1_q_net_x5;
  frame_pixel_2_at_offset_3 <= x12_bit_bin_value_2_q_net_x5;
  frame_pixel_3_at_offset_3 <= x12_bit_bin_value_3_q_net_x5;
  frame_pixel_4_at_offset_3 <= x12_bit_bin_value_4_q_net_x5;
  frame_pixel_5_at_offset_3 <= x12_bit_bin_value_5_q_net_x5;
  frame_pixel_6_at_offset_3 <= x12_bit_bin_value_6_q_net_x5;
  frame_pixel_7_at_offset_3 <= x12_bit_bin_value_7_q_net_x5;
  frame_pixel_8_at_offset_3 <= x12_bit_bin_value_8_q_net_x5;
  frame_pixel_9_at_offset_3 <= x12_bit_bin_value_9_q_net_x5;
  frame_pixel_10_at_offset_3 <= x12_bit_bin_value_10_q_net_x5;
  frame_pixel_11_at_offset_3 <= x12_bit_bin_value_11_q_net_x5;
  frame_pixel_0_at_offset_4 <= x12_bit_bin_value_0_q_net_x4;
  frame_pixel_1_at_offset_4 <= x12_bit_bin_value_1_q_net_x4;
  frame_pixel_2_at_offset_4 <= x12_bit_bin_value_2_q_net_x4;
  frame_pixel_3_at_offset_4 <= x12_bit_bin_value_3_q_net_x4;
  frame_pixel_4_at_offset_4 <= x12_bit_bin_value_4_q_net_x4;
  frame_pixel_5_at_offset_4 <= x12_bit_bin_value_5_q_net_x4;
  frame_pixel_6_at_offset_4 <= x12_bit_bin_value_6_q_net_x4;
  frame_pixel_7_at_offset_4 <= x12_bit_bin_value_7_q_net_x4;
  frame_pixel_8_at_offset_4 <= x12_bit_bin_value_8_q_net_x4;
  frame_pixel_9_at_offset_4 <= x12_bit_bin_value_9_q_net_x4;
  frame_pixel_10_at_offset_4 <= x12_bit_bin_value_10_q_net_x4;
  frame_pixel_11_at_offset_4 <= x12_bit_bin_value_11_q_net_x4;
  weight_0_at_offset_0 <= x12_bit_bin_value_0_q_net_x3;
  weight_1_at_offset_0 <= x12_bit_bin_value_1_q_net_x3;
  weight_2_at_offset_0 <= x12_bit_bin_value_2_q_net_x3;
  weight_3_at_offset_0 <= x12_bit_bin_value_3_q_net_x3;
  weight_4_at_offset_0 <= x12_bit_bin_value_4_q_net_x3;
  weight_5_at_offset_0 <= x12_bit_bin_value_5_q_net_x3;
  weight_6_at_offset_0 <= x12_bit_bin_value_6_q_net_x3;
  weight_7_at_offset_0 <= x12_bit_bin_value_7_q_net_x3;
  weight_8_at_offset_0 <= x12_bit_bin_value_8_q_net_x3;
  weight_9_at_offset_0 <= x12_bit_bin_value_9_q_net_x3;
  weight_10_at_offset_0 <= x12_bit_bin_value_10_q_net_x3;
  weight_11_at_offset_0 <= x12_bit_bin_value_11_q_net_x3;
  weight_0_at_offset_1 <= x12_bit_bin_value_0_q_net_x2;
  weight_1_at_offset_1 <= x12_bit_bin_value_1_q_net_x2;
  weight_2_at_offset_1 <= x12_bit_bin_value_2_q_net_x2;
  weight_3_at_offset_1 <= x12_bit_bin_value_3_q_net_x2;
  weight_4_at_offset_1 <= x12_bit_bin_value_4_q_net_x2;
  weight_5_at_offset_1 <= x12_bit_bin_value_5_q_net_x2;
  weight_6_at_offset_1 <= x12_bit_bin_value_6_q_net_x2;
  weight_7_at_offset_1 <= x12_bit_bin_value_7_q_net_x2;
  weight_8_at_offset_1 <= x12_bit_bin_value_8_q_net_x2;
  weight_9_at_offset_1 <= x12_bit_bin_value_9_q_net_x2;
  weight_10_at_offset_1 <= x12_bit_bin_value_10_q_net_x2;
  weight_11_at_offset_1 <= x12_bit_bin_value_11_q_net_x2;
  weight_0_at_offset_2 <= x12_bit_bin_value_0_q_net_x1;
  weight_1_at_offset_2 <= x12_bit_bin_value_1_q_net_x1;
  weight_2_at_offset_2 <= x12_bit_bin_value_2_q_net_x1;
  weight_3_at_offset_2 <= x12_bit_bin_value_3_q_net_x1;
  weight_4_at_offset_2 <= x12_bit_bin_value_4_q_net_x1;
  weight_5_at_offset_2 <= x12_bit_bin_value_5_q_net_x1;
  weight_6_at_offset_2 <= x12_bit_bin_value_6_q_net_x1;
  weight_7_at_offset_2 <= x12_bit_bin_value_7_q_net_x1;
  weight_8_at_offset_2 <= x12_bit_bin_value_8_q_net_x1;
  weight_9_at_offset_2 <= x12_bit_bin_value_9_q_net_x1;
  weight_10_at_offset_2 <= x12_bit_bin_value_10_q_net_x1;
  weight_11_at_offset_2 <= x12_bit_bin_value_11_q_net_x1;
  weight_0_at_offset_3 <= x12_bit_bin_value_0_q_net_x0;
  weight_1_at_offset_3 <= x12_bit_bin_value_1_q_net_x0;
  weight_2_at_offset_3 <= x12_bit_bin_value_2_q_net_x0;
  weight_3_at_offset_3 <= x12_bit_bin_value_3_q_net_x0;
  weight_4_at_offset_3 <= x12_bit_bin_value_4_q_net_x0;
  weight_5_at_offset_3 <= x12_bit_bin_value_5_q_net_x0;
  weight_6_at_offset_3 <= x12_bit_bin_value_6_q_net_x0;
  weight_7_at_offset_3 <= x12_bit_bin_value_7_q_net_x0;
  weight_8_at_offset_3 <= x12_bit_bin_value_8_q_net_x0;
  weight_9_at_offset_3 <= x12_bit_bin_value_9_q_net_x0;
  weight_10_at_offset_3 <= x12_bit_bin_value_10_q_net_x0;
  weight_11_at_offset_3 <= x12_bit_bin_value_11_q_net_x0;
  weight_0_at_offset_4 <= x12_bit_bin_value_0_q_net;
  weight_1_at_offset_4 <= x12_bit_bin_value_1_q_net;
  weight_2_at_offset_4 <= x12_bit_bin_value_2_q_net;
  weight_3_at_offset_4 <= x12_bit_bin_value_3_q_net;
  weight_4_at_offset_4 <= x12_bit_bin_value_4_q_net;
  weight_5_at_offset_4 <= x12_bit_bin_value_5_q_net;
  weight_6_at_offset_4 <= x12_bit_bin_value_6_q_net;
  weight_7_at_offset_4 <= x12_bit_bin_value_7_q_net;
  weight_8_at_offset_4 <= x12_bit_bin_value_8_q_net;
  weight_9_at_offset_4 <= x12_bit_bin_value_9_q_net;
  weight_10_at_offset_4 <= x12_bit_bin_value_10_q_net;
  weight_11_at_offset_4 <= x12_bit_bin_value_11_q_net;
  valid_data <= data_valid_out_delay_q_net;
  dual_port_ram_0_douta_net_x0 <= data_in_ram_0;
  dual_port_ram_1_douta_net_x0 <= data_in_ram_1;
  dual_port_ram_2_douta_net_x0 <= data_in_ram_2;
  dual_port_ram_3_douta_net_x0 <= data_in_ram_3;
  dual_port_ram_4_douta_net_x0 <= data_in_ram_4;
  convert_to_bool_dout_net <= frame_valid_in;
  dual_port_ram_0_douta_net <= kernel_data_in_ram_0;
  dual_port_ram_1_douta_net <= kernel_data_in_ram_1;
  dual_port_ram_2_douta_net <= kernel_data_in_ram_2;
  dual_port_ram_3_douta_net <= kernel_data_in_ram_3;
  dual_port_ram_4_douta_net <= kernel_data_in_ram_4;
  convert_to_bool_dout_net_x0 <= kernel_valid_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  frame_ram_slicer : entity xil_defaultlib.mh_frame_ram_slicer 
  port map (
    data_in_ram_0 => dual_port_ram_0_douta_net_x0,
    data_in_ram_1 => dual_port_ram_1_douta_net_x0,
    data_in_ram_2 => dual_port_ram_2_douta_net_x0,
    data_in_ram_3 => dual_port_ram_3_douta_net_x0,
    data_in_ram_4 => dual_port_ram_4_douta_net_x0,
    valid_in => convert_to_bool_dout_net,
    read_enable => read_out_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    frame_12_bit_bin_value_0_ram_0 => delay_5_q_net_x0,
    frame_12_bit_bin_value_1_ram_0 => delay_4_q_net_x0,
    frame_12_bit_bin_value_2_ram_0 => delay_3_q_net_x0,
    frame_12_bit_bin_value_3_ram_0 => delay_2_q_net_x0,
    frame_12_bit_bin_value_4_ram_0 => delay_1_q_net_x0,
    frame_12_bit_bin_value_5_ram_0 => delay_0_q_net_x0,
    frame_12_bit_bin_value_6_ram_0 => delay_11_q_net_x0,
    frame_12_bit_bin_value_7_ram_0 => delay_10_q_net_x0,
    frame_12_bit_bin_value_8_ram_0 => delay_9_q_net_x0,
    frame_12_bit_bin_value_9_ram_0 => delay_8_q_net_x0,
    frame_12_bit_bin_value_10_ram_0 => delay_7_q_net_x0,
    frame_12_bit_bin_value_11_ram_0 => delay_6_q_net_x0,
    frame_12_bit_bin_value_0_ram_1 => delay_19_q_net_x0,
    frame_12_bit_bin_value_1_ram_1 => delay_18_q_net_x0,
    frame_12_bit_bin_value_2_ram_1 => delay_17_q_net_x0,
    frame_12_bit_bin_value_3_ram_1 => delay_16_q_net_x0,
    frame_12_bit_bin_value_4_ram_1 => delay_13_q_net_x0,
    frame_12_bit_bin_value_5_ram_1 => delay_12_q_net_x0,
    frame_12_bit_bin_value_6_ram_1 => delay_15_q_net_x0,
    frame_12_bit_bin_value_7_ram_1 => delay_14_q_net_x0,
    frame_12_bit_bin_value_8_ram_1 => delay_23_q_net_x0,
    frame_12_bit_bin_value_9_ram_1 => delay_22_q_net_x0,
    frame_12_bit_bin_value_10_ram_1 => delay_21_q_net_x0,
    frame_12_bit_bin_value_11_ram_1 => delay_20_q_net_x0,
    frame_12_bit_bin_value_0_ram_2 => delay_43_q_net_x0,
    frame_12_bit_bin_value_1_ram_2 => delay_42_q_net_x0,
    frame_12_bit_bin_value_2_ram_2 => delay_41_q_net_x0,
    frame_12_bit_bin_value_3_ram_2 => delay_36_q_net_x0,
    frame_12_bit_bin_value_4_ram_2 => delay_25_q_net_x0,
    frame_12_bit_bin_value_5_ram_2 => delay_24_q_net_x0,
    frame_12_bit_bin_value_6_ram_2 => delay_27_q_net_x0,
    frame_12_bit_bin_value_7_ram_2 => delay_26_q_net_x0,
    frame_12_bit_bin_value_8_ram_2 => delay_47_q_net_x0,
    frame_12_bit_bin_value_9_ram_2 => delay_46_q_net_x0,
    frame_12_bit_bin_value_10_ram_2 => delay_45_q_net_x0,
    frame_12_bit_bin_value_11_ram_2 => delay_44_q_net_x0,
    frame_12_bit_bin_value_0_ram_3 => delay_35_q_net_x0,
    frame_12_bit_bin_value_1_ram_3 => delay_34_q_net_x0,
    frame_12_bit_bin_value_2_ram_3 => delay_33_q_net_x0,
    frame_12_bit_bin_value_3_ram_3 => delay_32_q_net_x0,
    frame_12_bit_bin_value_4_ram_3 => delay_29_q_net_x0,
    frame_12_bit_bin_value_5_ram_3 => delay_28_q_net_x0,
    frame_12_bit_bin_value_6_ram_3 => delay_31_q_net_x0,
    frame_12_bit_bin_value_7_ram_3 => delay_30_q_net_x0,
    frame_12_bit_bin_value_8_ram_3 => delay_40_q_net_x0,
    frame_12_bit_bin_value_9_ram_3 => delay_39_q_net_x0,
    frame_12_bit_bin_value_10_ram_3 => delay_38_q_net_x0,
    frame_12_bit_bin_value_11_ram_3 => delay_37_q_net_x0,
    frame_12_bit_bin_value_0_ram_4 => delay_67_q_net,
    frame_12_bit_bin_value_1_ram_4 => delay_66_q_net,
    frame_12_bit_bin_value_2_ram_4 => delay_65_q_net,
    frame_12_bit_bin_value_3_ram_4 => delay_60_q_net,
    frame_12_bit_bin_value_4_ram_4 => delay_49_q_net_x0,
    frame_12_bit_bin_value_5_ram_4 => delay_48_q_net_x0,
    frame_12_bit_bin_value_6_ram_4 => delay_51_q_net_x0,
    frame_12_bit_bin_value_7_ram_4 => delay_50_q_net_x0,
    frame_12_bit_bin_value_8_ram_4 => delay_71_q_net,
    frame_12_bit_bin_value_9_ram_4 => delay_70_q_net,
    frame_12_bit_bin_value_10_ram_4 => delay_69_q_net,
    frame_12_bit_bin_value_11_ram_4 => delay_68_q_net,
    valid_out => valid_sync_y_net_x0,
    wrote_to_last_fifo_ram_0 => logical_y_net_x8,
    wrote_to_last_fifo_ram_1 => logical_y_net_x7,
    wrote_to_last_fifo_ram_2 => logical_y_net_x6,
    wrote_to_last_fifo_ram_3 => logical_y_net_x5,
    wrote_to_last_fifo_ram_4 => logical_y_net_x4
  );
  kernel_ram_slicer : entity xil_defaultlib.mh_kernel_ram_slicer 
  port map (
    kernel_data_in_ram_0 => dual_port_ram_0_douta_net,
    kernel_data_in_ram_1 => dual_port_ram_1_douta_net,
    kernel_data_in_ram_2 => dual_port_ram_2_douta_net,
    kernel_data_in_ram_3 => dual_port_ram_3_douta_net,
    kernel_data_in_ram_4 => dual_port_ram_4_douta_net,
    valid_in => convert_to_bool_dout_net_x0,
    read_enable => read_out_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0_ram_0 => delay_3_q_net,
    kernel_18_bit_value_1_ram_0 => delay_2_q_net,
    kernel_18_bit_value_2_ram_0 => delay_1_q_net,
    kernel_18_bit_value_3_ram_0 => delay_0_q_net,
    kernel_18_bit_value_4_ram_0 => delay_7_q_net,
    kernel_18_bit_value_5_ram_0 => delay_6_q_net,
    kernel_18_bit_value_6_ram_0 => delay_5_q_net,
    kernel_18_bit_value_7_ram_0 => delay_4_q_net,
    kernel_18_bit_value_8_ram_0 => delay_11_q_net,
    kernel_18_bit_value_9_ram_0 => delay_10_q_net,
    kernel_18_bit_value_10_ram_0 => delay_9_q_net,
    kernel_18_bit_value_11_ram_0 => delay_8_q_net,
    kernel_18_bit_value_0_ram_1 => delay_17_q_net,
    kernel_18_bit_value_1_ram_1 => delay_16_q_net,
    kernel_18_bit_value_2_ram_1 => delay_13_q_net,
    kernel_18_bit_value_3_ram_1 => delay_12_q_net,
    kernel_18_bit_value_4_ram_1 => delay_21_q_net,
    kernel_18_bit_value_5_ram_1 => delay_20_q_net,
    kernel_18_bit_value_6_ram_1 => delay_19_q_net,
    kernel_18_bit_value_7_ram_1 => delay_18_q_net,
    kernel_18_bit_value_8_ram_1 => delay_15_q_net,
    kernel_18_bit_value_9_ram_1 => delay_14_q_net,
    kernel_18_bit_value_10_ram_1 => delay_23_q_net,
    kernel_18_bit_value_11_ram_1 => delay_22_q_net,
    kernel_18_bit_value_0_ram_2 => delay_29_q_net,
    kernel_18_bit_value_1_ram_2 => delay_28_q_net,
    kernel_18_bit_value_2_ram_2 => delay_25_q_net,
    kernel_18_bit_value_3_ram_2 => delay_24_q_net,
    kernel_18_bit_value_4_ram_2 => delay_33_q_net,
    kernel_18_bit_value_5_ram_2 => delay_32_q_net,
    kernel_18_bit_value_6_ram_2 => delay_31_q_net,
    kernel_18_bit_value_7_ram_2 => delay_30_q_net,
    kernel_18_bit_value_8_ram_2 => delay_27_q_net,
    kernel_18_bit_value_9_ram_2 => delay_26_q_net,
    kernel_18_bit_value_10_ram_2 => delay_35_q_net,
    kernel_18_bit_value_11_ram_2 => delay_34_q_net,
    kernel_18_bit_value_0_ram_3 => delay_41_q_net,
    kernel_18_bit_value_1_ram_3 => delay_40_q_net,
    kernel_18_bit_value_2_ram_3 => delay_37_q_net,
    kernel_18_bit_value_3_ram_3 => delay_36_q_net,
    kernel_18_bit_value_4_ram_3 => delay_45_q_net,
    kernel_18_bit_value_5_ram_3 => delay_44_q_net,
    kernel_18_bit_value_6_ram_3 => delay_43_q_net,
    kernel_18_bit_value_7_ram_3 => delay_42_q_net,
    kernel_18_bit_value_8_ram_3 => delay_39_q_net,
    kernel_18_bit_value_9_ram_3 => delay_38_q_net,
    kernel_18_bit_value_10_ram_3 => delay_47_q_net,
    kernel_18_bit_value_11_ram_3 => delay_46_q_net,
    kernel_18_bit_value_0_ram_4 => delay_53_q_net,
    kernel_18_bit_value_1_ram_4 => delay_52_q_net,
    kernel_18_bit_value_2_ram_4 => delay_49_q_net,
    kernel_18_bit_value_3_ram_4 => delay_48_q_net,
    kernel_18_bit_value_4_ram_4 => delay_57_q_net,
    kernel_18_bit_value_5_ram_4 => delay_56_q_net,
    kernel_18_bit_value_6_ram_4 => delay_55_q_net,
    kernel_18_bit_value_7_ram_4 => delay_54_q_net,
    kernel_18_bit_value_8_ram_4 => delay_51_q_net,
    kernel_18_bit_value_9_ram_4 => delay_50_q_net,
    kernel_18_bit_value_10_ram_4 => delay_59_q_net,
    kernel_18_bit_value_11_ram_4 => delay_58_q_net,
    valid_out => valid_sync_y_net,
    wrote_to_last_fifo_ram_0 => logical_y_net_x3,
    wrote_to_last_fifo_ram_1 => logical_y_net_x2,
    wrote_to_last_fifo_ram_2 => logical_y_net_x1,
    wrote_to_last_fifo_ram_3 => logical_y_net_x0,
    wrote_to_last_fifo_ram_4 => logical_y_net,
    wrote_to_last_fifo_trigger => last_fifo_written_to_1_q_net
  );
  subsystem1 : entity xil_defaultlib.mh_subsystem1 
  port map (
    frame_12_bit_bin_value_0 => delay_5_q_net_x0,
    frame_12_bit_bin_value_1 => delay_4_q_net_x0,
    frame_12_bit_bin_value_2 => delay_3_q_net_x0,
    frame_12_bit_bin_value_3 => delay_2_q_net_x0,
    frame_12_bit_bin_value_4 => delay_1_q_net_x0,
    frame_12_bit_bin_value_5 => delay_0_q_net_x0,
    frame_12_bit_bin_value_6 => delay_11_q_net_x0,
    frame_12_bit_bin_value_7 => delay_10_q_net_x0,
    frame_12_bit_bin_value_8 => delay_9_q_net_x0,
    frame_12_bit_bin_value_9 => delay_8_q_net_x0,
    frame_12_bit_bin_value_10 => delay_7_q_net_x0,
    frame_12_bit_bin_value_11 => delay_6_q_net_x0,
    frame_12_bit_bin_value_12 => delay_19_q_net_x0,
    frame_12_bit_bin_value_13 => delay_18_q_net_x0,
    frame_12_bit_bin_value_14 => delay_17_q_net_x0,
    frame_12_bit_bin_value_15 => delay_16_q_net_x0,
    frame_12_bit_bin_value_16 => delay_13_q_net_x0,
    frame_12_bit_bin_value_17 => delay_12_q_net_x0,
    frame_12_bit_bin_value_18 => delay_15_q_net_x0,
    frame_12_bit_bin_value_19 => delay_14_q_net_x0,
    frame_12_bit_bin_value_20 => delay_23_q_net_x0,
    frame_12_bit_bin_value_21 => delay_22_q_net_x0,
    frame_12_bit_bin_value_22 => delay_21_q_net_x0,
    frame_12_bit_bin_value_23 => delay_20_q_net_x0,
    frame_12_bit_bin_value_24 => delay_43_q_net_x0,
    frame_12_bit_bin_value_25 => delay_42_q_net_x0,
    frame_12_bit_bin_value_26 => delay_41_q_net_x0,
    frame_12_bit_bin_value_27 => delay_36_q_net_x0,
    frame_12_bit_bin_value_28 => delay_25_q_net_x0,
    frame_12_bit_bin_value_29 => delay_24_q_net_x0,
    frame_12_bit_bin_value_30 => delay_27_q_net_x0,
    frame_12_bit_bin_value_31 => delay_26_q_net_x0,
    frame_12_bit_bin_value_32 => delay_47_q_net_x0,
    frame_12_bit_bin_value_33 => delay_46_q_net_x0,
    frame_12_bit_bin_value_34 => delay_45_q_net_x0,
    frame_12_bit_bin_value_35 => delay_44_q_net_x0,
    frame_12_bit_bin_value_36 => delay_35_q_net_x0,
    frame_12_bit_bin_value_37 => delay_34_q_net_x0,
    frame_12_bit_bin_value_38 => delay_33_q_net_x0,
    frame_12_bit_bin_value_39 => delay_32_q_net_x0,
    frame_12_bit_bin_value_40 => delay_29_q_net_x0,
    frame_12_bit_bin_value_41 => delay_28_q_net_x0,
    frame_12_bit_bin_value_42 => delay_31_q_net_x0,
    frame_12_bit_bin_value_43 => delay_30_q_net_x0,
    frame_12_bit_bin_value_44 => delay_40_q_net_x0,
    frame_12_bit_bin_value_45 => delay_39_q_net_x0,
    frame_12_bit_bin_value_46 => delay_38_q_net_x0,
    frame_12_bit_bin_value_47 => delay_37_q_net_x0,
    frame_12_bit_bin_value_48 => delay_67_q_net,
    frame_12_bit_bin_value_49 => delay_66_q_net,
    frame_12_bit_bin_value_50 => delay_65_q_net,
    frame_12_bit_bin_value_51 => delay_60_q_net,
    frame_12_bit_bin_value_52 => delay_49_q_net_x0,
    frame_12_bit_bin_value_53 => delay_48_q_net_x0,
    frame_12_bit_bin_value_54 => delay_51_q_net_x0,
    frame_12_bit_bin_value_55 => delay_50_q_net_x0,
    frame_12_bit_bin_value_56 => delay_71_q_net,
    frame_12_bit_bin_value_57 => delay_70_q_net,
    frame_12_bit_bin_value_58 => delay_69_q_net,
    frame_12_bit_bin_value_59 => delay_68_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    frame_12_bit_value_0 => x12_bit_bin_value_0_q_net_x8,
    frame_12_bit_value_1 => x12_bit_bin_value_1_q_net_x8,
    frame_12_bit_value_2 => x12_bit_bin_value_2_q_net_x8,
    frame_12_bit_value_3 => x12_bit_bin_value_3_q_net_x8,
    frame_12_bit_value_4 => x12_bit_bin_value_4_q_net_x8,
    frame_12_bit_value_5 => x12_bit_bin_value_5_q_net_x8,
    frame_12_bit_value_6 => x12_bit_bin_value_6_q_net_x8,
    frame_12_bit_value_7 => x12_bit_bin_value_7_q_net_x8,
    frame_12_bit_value_8 => x12_bit_bin_value_8_q_net_x8,
    frame_12_bit_value_9 => x12_bit_bin_value_9_q_net_x8,
    frame_12_bit_value_10 => x12_bit_bin_value_10_q_net_x8,
    frame_12_bit_value_11 => x12_bit_bin_value_11_q_net_x8,
    frame_12_bit_value_12 => x12_bit_bin_value_0_q_net_x7,
    frame_12_bit_value_13 => x12_bit_bin_value_1_q_net_x7,
    frame_12_bit_value_14 => x12_bit_bin_value_2_q_net_x7,
    frame_12_bit_value_15 => x12_bit_bin_value_3_q_net_x7,
    frame_12_bit_value_16 => x12_bit_bin_value_4_q_net_x7,
    frame_12_bit_value_17 => x12_bit_bin_value_5_q_net_x7,
    frame_12_bit_value_18 => x12_bit_bin_value_6_q_net_x7,
    frame_12_bit_value_19 => x12_bit_bin_value_7_q_net_x7,
    frame_12_bit_value_20 => x12_bit_bin_value_8_q_net_x7,
    frame_12_bit_value_21 => x12_bit_bin_value_9_q_net_x7,
    frame_12_bit_value_22 => x12_bit_bin_value_10_q_net_x7,
    frame_12_bit_value_23 => x12_bit_bin_value_11_q_net_x7,
    frame_12_bit_value_24 => x12_bit_bin_value_0_q_net_x6,
    frame_12_bit_value_25 => x12_bit_bin_value_1_q_net_x6,
    frame_12_bit_value_26 => x12_bit_bin_value_2_q_net_x6,
    frame_12_bit_value_27 => x12_bit_bin_value_3_q_net_x6,
    frame_12_bit_value_28 => x12_bit_bin_value_4_q_net_x6,
    frame_12_bit_value_29 => x12_bit_bin_value_5_q_net_x6,
    frame_12_bit_value_30 => x12_bit_bin_value_6_q_net_x6,
    frame_12_bit_value_31 => x12_bit_bin_value_7_q_net_x6,
    frame_12_bit_value_32 => x12_bit_bin_value_8_q_net_x6,
    frame_12_bit_value_33 => x12_bit_bin_value_9_q_net_x6,
    frame_12_bit_value_34 => x12_bit_bin_value_10_q_net_x6,
    frame_12_bit_value_35 => x12_bit_bin_value_11_q_net_x6,
    frame_12_bit_value_36 => x12_bit_bin_value_0_q_net_x5,
    frame_12_bit_value_37 => x12_bit_bin_value_1_q_net_x5,
    frame_12_bit_value_38 => x12_bit_bin_value_2_q_net_x5,
    frame_12_bit_value_39 => x12_bit_bin_value_3_q_net_x5,
    frame_12_bit_value_40 => x12_bit_bin_value_4_q_net_x5,
    frame_12_bit_value_41 => x12_bit_bin_value_5_q_net_x5,
    frame_12_bit_value_42 => x12_bit_bin_value_6_q_net_x5,
    frame_12_bit_value_43 => x12_bit_bin_value_7_q_net_x5,
    frame_12_bit_value_44 => x12_bit_bin_value_8_q_net_x5,
    frame_12_bit_value_45 => x12_bit_bin_value_9_q_net_x5,
    frame_12_bit_value_46 => x12_bit_bin_value_10_q_net_x5,
    frame_12_bit_value_47 => x12_bit_bin_value_11_q_net_x5,
    frame_12_bit_value_48 => x12_bit_bin_value_0_q_net_x4,
    frame_12_bit_value_49 => x12_bit_bin_value_1_q_net_x4,
    frame_12_bit_value_50 => x12_bit_bin_value_2_q_net_x4,
    frame_12_bit_value_51 => x12_bit_bin_value_3_q_net_x4,
    frame_12_bit_value_52 => x12_bit_bin_value_4_q_net_x4,
    frame_12_bit_value_53 => x12_bit_bin_value_5_q_net_x4,
    frame_12_bit_value_54 => x12_bit_bin_value_6_q_net_x4,
    frame_12_bit_value_55 => x12_bit_bin_value_7_q_net_x4,
    frame_12_bit_value_56 => x12_bit_bin_value_8_q_net_x4,
    frame_12_bit_value_57 => x12_bit_bin_value_9_q_net_x4,
    frame_12_bit_value_58 => x12_bit_bin_value_10_q_net_x4,
    frame_12_bit_value_59 => x12_bit_bin_value_11_q_net_x4
  );
  subsystem2 : entity xil_defaultlib.mh_subsystem2 
  port map (
    kernel_18_bit_bin_value_0 => delay_3_q_net,
    kernel_18_bit_bin_value_1 => delay_2_q_net,
    kernel_18_bit_bin_value_2 => delay_1_q_net,
    kernel_18_bit_bin_value_3 => delay_0_q_net,
    kernel_18_bit_bin_value_4 => delay_7_q_net,
    kernel_18_bit_bin_value_5 => delay_6_q_net,
    kernel_18_bit_bin_value_6 => delay_5_q_net,
    kernel_18_bit_bin_value_7 => delay_4_q_net,
    kernel_18_bit_bin_value_8 => delay_11_q_net,
    kernel_18_bit_bin_value_9 => delay_10_q_net,
    kernel_18_bit_bin_value_10 => delay_9_q_net,
    kernel_18_bit_bin_value_11 => delay_8_q_net,
    kernel_18_bit_bin_value_12 => delay_17_q_net,
    kernel_18_bit_bin_value_13 => delay_16_q_net,
    kernel_18_bit_bin_value_14 => delay_13_q_net,
    kernel_18_bit_bin_value_15 => delay_12_q_net,
    kernel_18_bit_bin_value_16 => delay_21_q_net,
    kernel_18_bit_bin_value_17 => delay_20_q_net,
    kernel_18_bit_bin_value_18 => delay_19_q_net,
    kernel_18_bit_bin_value_19 => delay_18_q_net,
    kernel_18_bit_bin_value_20 => delay_15_q_net,
    kernel_18_bit_bin_value_21 => delay_14_q_net,
    kernel_18_bit_bin_value_22 => delay_23_q_net,
    kernel_18_bit_bin_value_23 => delay_22_q_net,
    kernel_18_bit_bin_value_24 => delay_29_q_net,
    kernel_18_bit_bin_value_25 => delay_28_q_net,
    kernel_18_bit_bin_value_26 => delay_25_q_net,
    kernel_18_bit_bin_value_27 => delay_24_q_net,
    kernel_18_bit_bin_value_28 => delay_33_q_net,
    kernel_18_bit_bin_value_29 => delay_32_q_net,
    kernel_18_bit_bin_value_30 => delay_31_q_net,
    kernel_18_bit_bin_value_31 => delay_30_q_net,
    kernel_18_bit_bin_value_32 => delay_27_q_net,
    kernel_18_bit_bin_value_33 => delay_26_q_net,
    kernel_18_bit_bin_value_34 => delay_35_q_net,
    kernel_18_bit_bin_value_35 => delay_34_q_net,
    kernel_18_bit_bin_value_36 => delay_41_q_net,
    kernel_18_bit_bin_value_37 => delay_40_q_net,
    kernel_18_bit_bin_value_38 => delay_37_q_net,
    kernel_18_bit_bin_value_39 => delay_36_q_net,
    kernel_18_bit_bin_value_40 => delay_45_q_net,
    kernel_18_bit_bin_value_41 => delay_44_q_net,
    kernel_18_bit_bin_value_42 => delay_43_q_net,
    kernel_18_bit_bin_value_43 => delay_42_q_net,
    kernel_18_bit_bin_value_44 => delay_39_q_net,
    kernel_18_bit_bin_value_45 => delay_38_q_net,
    kernel_18_bit_bin_value_46 => delay_47_q_net,
    kernel_18_bit_bin_value_47 => delay_46_q_net,
    kernel_18_bit_bin_value_48 => delay_53_q_net,
    kernel_18_bit_bin_value_49 => delay_52_q_net,
    kernel_18_bit_bin_value_50 => delay_49_q_net,
    kernel_18_bit_bin_value_51 => delay_48_q_net,
    kernel_18_bit_bin_value_52 => delay_57_q_net,
    kernel_18_bit_bin_value_53 => delay_56_q_net,
    kernel_18_bit_bin_value_54 => delay_55_q_net,
    kernel_18_bit_bin_value_55 => delay_54_q_net,
    kernel_18_bit_bin_value_56 => delay_51_q_net,
    kernel_18_bit_bin_value_57 => delay_50_q_net,
    kernel_18_bit_bin_value_58 => delay_59_q_net,
    kernel_18_bit_bin_value_59 => delay_58_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_18_bit_value_0 => x12_bit_bin_value_0_q_net_x3,
    kernel_18_bit_value_1 => x12_bit_bin_value_1_q_net_x3,
    kernel_18_bit_value_2 => x12_bit_bin_value_2_q_net_x3,
    kernel_18_bit_value_3 => x12_bit_bin_value_3_q_net_x3,
    kernel_18_bit_value_4 => x12_bit_bin_value_4_q_net_x3,
    kernel_18_bit_value_5 => x12_bit_bin_value_5_q_net_x3,
    kernel_18_bit_value_6 => x12_bit_bin_value_6_q_net_x3,
    kernel_18_bit_value_7 => x12_bit_bin_value_7_q_net_x3,
    kernel_18_bit_value_8 => x12_bit_bin_value_8_q_net_x3,
    kernel_18_bit_value_9 => x12_bit_bin_value_9_q_net_x3,
    kernel_18_bit_value_10 => x12_bit_bin_value_10_q_net_x3,
    kernel_18_bit_value_11 => x12_bit_bin_value_11_q_net_x3,
    kernel_18_bit_value_12 => x12_bit_bin_value_0_q_net_x2,
    kernel_18_bit_value_13 => x12_bit_bin_value_1_q_net_x2,
    kernel_18_bit_value_14 => x12_bit_bin_value_2_q_net_x2,
    kernel_18_bit_value_15 => x12_bit_bin_value_3_q_net_x2,
    kernel_18_bit_value_16 => x12_bit_bin_value_4_q_net_x2,
    kernel_18_bit_value_17 => x12_bit_bin_value_5_q_net_x2,
    kernel_18_bit_value_18 => x12_bit_bin_value_6_q_net_x2,
    kernel_18_bit_value_19 => x12_bit_bin_value_7_q_net_x2,
    kernel_18_bit_value_20 => x12_bit_bin_value_8_q_net_x2,
    kernel_18_bit_value_21 => x12_bit_bin_value_9_q_net_x2,
    kernel_18_bit_value_22 => x12_bit_bin_value_10_q_net_x2,
    kernel_18_bit_value_23 => x12_bit_bin_value_11_q_net_x2,
    kernel_18_bit_value_24 => x12_bit_bin_value_0_q_net_x1,
    kernel_18_bit_value_25 => x12_bit_bin_value_1_q_net_x1,
    kernel_18_bit_value_26 => x12_bit_bin_value_2_q_net_x1,
    kernel_18_bit_value_27 => x12_bit_bin_value_3_q_net_x1,
    kernel_18_bit_value_28 => x12_bit_bin_value_4_q_net_x1,
    kernel_18_bit_value_29 => x12_bit_bin_value_5_q_net_x1,
    kernel_18_bit_value_30 => x12_bit_bin_value_6_q_net_x1,
    kernel_18_bit_value_31 => x12_bit_bin_value_7_q_net_x1,
    kernel_18_bit_value_32 => x12_bit_bin_value_8_q_net_x1,
    kernel_18_bit_value_33 => x12_bit_bin_value_9_q_net_x1,
    kernel_18_bit_value_34 => x12_bit_bin_value_10_q_net_x1,
    kernel_18_bit_value_35 => x12_bit_bin_value_11_q_net_x1,
    kernel_18_bit_value_36 => x12_bit_bin_value_0_q_net_x0,
    kernel_18_bit_value_37 => x12_bit_bin_value_1_q_net_x0,
    kernel_18_bit_value_38 => x12_bit_bin_value_2_q_net_x0,
    kernel_18_bit_value_39 => x12_bit_bin_value_3_q_net_x0,
    kernel_18_bit_value_40 => x12_bit_bin_value_4_q_net_x0,
    kernel_18_bit_value_41 => x12_bit_bin_value_5_q_net_x0,
    kernel_18_bit_value_42 => x12_bit_bin_value_6_q_net_x0,
    kernel_18_bit_value_43 => x12_bit_bin_value_7_q_net_x0,
    kernel_18_bit_value_44 => x12_bit_bin_value_8_q_net_x0,
    kernel_18_bit_value_45 => x12_bit_bin_value_9_q_net_x0,
    kernel_18_bit_value_46 => x12_bit_bin_value_10_q_net_x0,
    kernel_18_bit_value_47 => x12_bit_bin_value_11_q_net_x0,
    kernel_18_bit_value_48 => x12_bit_bin_value_0_q_net,
    kernel_18_bit_value_49 => x12_bit_bin_value_1_q_net,
    kernel_18_bit_value_50 => x12_bit_bin_value_2_q_net,
    kernel_18_bit_value_51 => x12_bit_bin_value_3_q_net,
    kernel_18_bit_value_52 => x12_bit_bin_value_4_q_net,
    kernel_18_bit_value_53 => x12_bit_bin_value_5_q_net,
    kernel_18_bit_value_54 => x12_bit_bin_value_6_q_net,
    kernel_18_bit_value_55 => x12_bit_bin_value_7_q_net,
    kernel_18_bit_value_56 => x12_bit_bin_value_8_q_net,
    kernel_18_bit_value_57 => x12_bit_bin_value_9_q_net,
    kernel_18_bit_value_58 => x12_bit_bin_value_10_q_net,
    kernel_18_bit_value_59 => x12_bit_bin_value_11_q_net
  );
  data_valid_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_out_y_net,
    clk => clk_net,
    ce => ce_net,
    q => data_valid_out_delay_q_net
  );
  read_out : entity xil_defaultlib.sysgen_logical_e0b850d218 
  port map (
    clr => '0',
    d0 => logical_y_net_x8,
    d1 => logical_y_net_x7,
    d2 => logical_y_net_x6,
    d3 => logical_y_net_x5,
    d4 => logical_y_net_x4,
    d5 => logical_y_net_x3,
    d6 => logical_y_net_x2,
    d7 => logical_y_net_x1,
    d8 => logical_y_net_x0,
    d9 => logical_y_net,
    d10 => last_fifo_written_to_1_q_net,
    clk => clk_net,
    ce => ce_net,
    y => read_out_y_net
  );
  valid_out : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => valid_sync_y_net_x0,
    d1 => valid_sync_y_net,
    clk => clk_net,
    ce => ce_net,
    y => valid_out_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_0 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    force_off : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_0;
architecture structural of mh_result_muxer_0 is 
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_0_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  last_kernel_op_net <= force_off;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  force_off_mux : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => last_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_1 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_1;
architecture structural of mh_result_muxer_1 is 
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_1_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_2 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_2;
architecture structural of mh_result_muxer_2 is 
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_1_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_3 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_3;
architecture structural of mh_result_muxer_3 is 
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_1_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_4 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_4;
architecture structural of mh_result_muxer_4 is 
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_1_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_5 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    force_off : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_5;
architecture structural of mh_result_muxer_5 is 
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal first_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux_y_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_1_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  first_kernel_op_net <= force_off;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  force_off_mux : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => first_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_6 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    force_off : in std_logic_vector( 1-1 downto 0 );
    force_off_2 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_6;
architecture structural of mh_result_muxer_6 is 
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal first_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux1_y_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_0_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  first_kernel_op_net <= force_off;
  last_kernel_op_net <= force_off_2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  force_off_mux : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => first_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux_y_net
  );
  force_off_mux1 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => last_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_7 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    force_off : in std_logic_vector( 1-1 downto 0 );
    force_off_2 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_7;
architecture structural of mh_result_muxer_7 is 
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal first_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux_y_net : std_logic_vector( 1-1 downto 0 );
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux1_y_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_0_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  first_kernel_op_net <= force_off;
  last_kernel_op_net <= force_off_2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  force_off_mux : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => first_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux_y_net
  );
  force_off_mux1 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => last_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 8
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_8 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    force_off : in std_logic_vector( 1-1 downto 0 );
    force_off_2 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_8;
architecture structural of mh_result_muxer_8 is 
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux1_y_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal force_off_mux_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal first_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_0_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  first_kernel_op_net <= force_off;
  last_kernel_op_net <= force_off_2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  force_off_mux : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => first_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux_y_net
  );
  force_off_mux1 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => last_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1/Result Muxer 9
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_result_muxer_9 is
  port (
    select_x0 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    force_off : in std_logic_vector( 1-1 downto 0 );
    force_off_2 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_slice_0_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_1_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_2_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_3_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_slice_4_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_result_muxer_9;
architecture structural of mh_result_muxer_9 is 
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal first_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal on_op_net : std_logic_vector( 1-1 downto 0 );
  signal off_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_valid_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux1_y_net : std_logic_vector( 1-1 downto 0 );
  signal force_off_mux_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_result_slice_0_valid <= enable_passthrough_case_1_y_net;
  kernel_result_slice_1_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_2_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_3_valid <= enable_passthrough_case_0_y_net;
  kernel_result_slice_4_valid <= enable_passthrough_case_0_y_net;
  disable_q_net <= select_x0;
  valid_data_delay_4_q_net <= valid;
  first_kernel_op_net <= force_off;
  last_kernel_op_net <= force_off_2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  case_0 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_0_y_net
  );
  case_1 : entity xil_defaultlib.sysgen_mux_ec1a7626fa 
  port map (
    clr => '0',
    sel => disable_q_net,
    d0 => off_op_net,
    d1 => on_op_net,
    clk => clk_net,
    ce => ce_net,
    y => case_1_y_net
  );
  delay_valid_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_valid_0_q_net
  );
  enable_passthrough_case_0 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_0_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_0_y_net
  );
  enable_passthrough_case_1 : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => case_1_y_net,
    d1 => delay_valid_0_q_net,
    d2 => force_off_mux_y_net,
    d3 => force_off_mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_passthrough_case_1_y_net
  );
  force_off_mux : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => first_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux_y_net
  );
  force_off_mux1 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => last_kernel_op_net,
    d0 => on_op_net,
    d1 => off_op_net,
    clk => clk_net,
    ce => ce_net,
    y => force_off_mux1_y_net
  );
  off : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => off_op_net
  );
  on_x0 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => on_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer/Determine Calculations Delay 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_determine_calculations_delay_1 is
  port (
    valid_data_in : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_valid_out_0_kernel_result_0 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_0 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_0 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_0 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_0 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_1 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_1 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_1 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_1 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_1 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_2 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_2 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_2 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_2 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_2 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_3 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_3 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_3 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_3 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_3 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_4 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_4 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_4 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_4 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_4 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_5 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_5 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_5 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_5 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_5 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_6 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_6 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_6 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_6 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_6 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_7 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_7 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_7 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_7 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_7 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_8 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_8 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_8 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_8 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_8 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_9 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_1_kernel_result_9 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_2_kernel_result_9 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_3_kernel_result_9 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_4_kernel_result_9 : out std_logic_vector( 1-1 downto 0 );
    slice_valid_out_0_kernel_result_10 : out std_logic_vector( 1-1 downto 0 )
  );
end mh_determine_calculations_delay_1;
architecture structural of mh_determine_calculations_delay_1 is 
  signal enable_passthrough_case_1_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_6_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_valid_out_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal enable_disable_kernels_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal logical3_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 10-1 downto 0 );
  signal valid_data_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_10_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal last_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_op_net : std_logic_vector( 10-1 downto 0 );
  signal disable_q_net : std_logic_vector( 1-1 downto 0 );
  signal first_kernel_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_row_enable_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal what_kernel_position_op_net : std_logic_vector( 12-1 downto 0 );
  signal valid_data_delay_11_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_kernel_op_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical2_y_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_5_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_7_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_3_q_net : std_logic_vector( 1-1 downto 0 );
  signal valid_data_delay_9_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_valid_out_0_kernel_result_0 <= enable_passthrough_case_0_y_net_x7;
  slice_valid_out_1_kernel_result_0 <= enable_passthrough_case_0_y_net_x7;
  slice_valid_out_2_kernel_result_0 <= enable_passthrough_case_0_y_net_x7;
  slice_valid_out_3_kernel_result_0 <= enable_passthrough_case_0_y_net_x7;
  slice_valid_out_4_kernel_result_0 <= enable_passthrough_case_0_y_net_x7;
  slice_valid_out_0_kernel_result_1 <= enable_passthrough_case_0_y_net_x6;
  slice_valid_out_1_kernel_result_1 <= enable_passthrough_case_0_y_net_x6;
  slice_valid_out_2_kernel_result_1 <= enable_passthrough_case_0_y_net_x6;
  slice_valid_out_3_kernel_result_1 <= enable_passthrough_case_0_y_net_x6;
  slice_valid_out_4_kernel_result_1 <= enable_passthrough_case_1_y_net_x7;
  slice_valid_out_0_kernel_result_2 <= enable_passthrough_case_0_y_net_x5;
  slice_valid_out_1_kernel_result_2 <= enable_passthrough_case_0_y_net_x5;
  slice_valid_out_2_kernel_result_2 <= enable_passthrough_case_0_y_net_x5;
  slice_valid_out_3_kernel_result_2 <= enable_passthrough_case_1_y_net_x6;
  slice_valid_out_4_kernel_result_2 <= enable_passthrough_case_1_y_net_x6;
  slice_valid_out_0_kernel_result_3 <= enable_passthrough_case_0_y_net_x4;
  slice_valid_out_1_kernel_result_3 <= enable_passthrough_case_0_y_net_x4;
  slice_valid_out_2_kernel_result_3 <= enable_passthrough_case_1_y_net_x5;
  slice_valid_out_3_kernel_result_3 <= enable_passthrough_case_1_y_net_x5;
  slice_valid_out_4_kernel_result_3 <= enable_passthrough_case_1_y_net_x5;
  slice_valid_out_0_kernel_result_4 <= enable_passthrough_case_0_y_net_x3;
  slice_valid_out_1_kernel_result_4 <= enable_passthrough_case_1_y_net_x4;
  slice_valid_out_2_kernel_result_4 <= enable_passthrough_case_1_y_net_x4;
  slice_valid_out_3_kernel_result_4 <= enable_passthrough_case_1_y_net_x4;
  slice_valid_out_4_kernel_result_4 <= enable_passthrough_case_1_y_net_x4;
  slice_valid_out_0_kernel_result_5 <= enable_passthrough_case_1_y_net_x3;
  slice_valid_out_1_kernel_result_5 <= enable_passthrough_case_1_y_net_x3;
  slice_valid_out_2_kernel_result_5 <= enable_passthrough_case_1_y_net_x3;
  slice_valid_out_3_kernel_result_5 <= enable_passthrough_case_1_y_net_x3;
  slice_valid_out_4_kernel_result_5 <= enable_passthrough_case_1_y_net_x3;
  slice_valid_out_0_kernel_result_6 <= enable_passthrough_case_1_y_net_x2;
  slice_valid_out_1_kernel_result_6 <= enable_passthrough_case_1_y_net_x2;
  slice_valid_out_2_kernel_result_6 <= enable_passthrough_case_1_y_net_x2;
  slice_valid_out_3_kernel_result_6 <= enable_passthrough_case_1_y_net_x2;
  slice_valid_out_4_kernel_result_6 <= enable_passthrough_case_0_y_net_x2;
  slice_valid_out_0_kernel_result_7 <= enable_passthrough_case_1_y_net_x1;
  slice_valid_out_1_kernel_result_7 <= enable_passthrough_case_1_y_net_x1;
  slice_valid_out_2_kernel_result_7 <= enable_passthrough_case_1_y_net_x1;
  slice_valid_out_3_kernel_result_7 <= enable_passthrough_case_0_y_net_x0;
  slice_valid_out_4_kernel_result_7 <= enable_passthrough_case_0_y_net_x0;
  slice_valid_out_0_kernel_result_8 <= enable_passthrough_case_1_y_net;
  slice_valid_out_1_kernel_result_8 <= enable_passthrough_case_1_y_net;
  slice_valid_out_2_kernel_result_8 <= enable_passthrough_case_0_y_net_x1;
  slice_valid_out_3_kernel_result_8 <= enable_passthrough_case_0_y_net_x1;
  slice_valid_out_4_kernel_result_8 <= enable_passthrough_case_0_y_net_x1;
  slice_valid_out_0_kernel_result_9 <= enable_passthrough_case_1_y_net_x0;
  slice_valid_out_1_kernel_result_9 <= enable_passthrough_case_0_y_net;
  slice_valid_out_2_kernel_result_9 <= enable_passthrough_case_0_y_net;
  slice_valid_out_3_kernel_result_9 <= enable_passthrough_case_0_y_net;
  slice_valid_out_4_kernel_result_9 <= enable_passthrough_case_0_y_net;
  slice_valid_out_0_kernel_result_10 <= last_out_q_net;
  data_valid_out_delay_q_net <= valid_data_in;
  switch_to_zero_y_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  result_muxer_0 : entity xil_defaultlib.mh_result_muxer_0 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    force_off => last_kernel_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_0_y_net_x7,
    kernel_result_slice_1_valid => enable_passthrough_case_0_y_net_x7,
    kernel_result_slice_2_valid => enable_passthrough_case_0_y_net_x7,
    kernel_result_slice_3_valid => enable_passthrough_case_0_y_net_x7,
    kernel_result_slice_4_valid => enable_passthrough_case_0_y_net_x7
  );
  result_muxer_1 : entity xil_defaultlib.mh_result_muxer_1 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_0_y_net_x6,
    kernel_result_slice_1_valid => enable_passthrough_case_0_y_net_x6,
    kernel_result_slice_2_valid => enable_passthrough_case_0_y_net_x6,
    kernel_result_slice_3_valid => enable_passthrough_case_0_y_net_x6,
    kernel_result_slice_4_valid => enable_passthrough_case_1_y_net_x7
  );
  result_muxer_2 : entity xil_defaultlib.mh_result_muxer_2 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_0_y_net_x5,
    kernel_result_slice_1_valid => enable_passthrough_case_0_y_net_x5,
    kernel_result_slice_2_valid => enable_passthrough_case_0_y_net_x5,
    kernel_result_slice_3_valid => enable_passthrough_case_1_y_net_x6,
    kernel_result_slice_4_valid => enable_passthrough_case_1_y_net_x6
  );
  result_muxer_3 : entity xil_defaultlib.mh_result_muxer_3 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_0_y_net_x4,
    kernel_result_slice_1_valid => enable_passthrough_case_0_y_net_x4,
    kernel_result_slice_2_valid => enable_passthrough_case_1_y_net_x5,
    kernel_result_slice_3_valid => enable_passthrough_case_1_y_net_x5,
    kernel_result_slice_4_valid => enable_passthrough_case_1_y_net_x5
  );
  result_muxer_4 : entity xil_defaultlib.mh_result_muxer_4 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_0_y_net_x3,
    kernel_result_slice_1_valid => enable_passthrough_case_1_y_net_x4,
    kernel_result_slice_2_valid => enable_passthrough_case_1_y_net_x4,
    kernel_result_slice_3_valid => enable_passthrough_case_1_y_net_x4,
    kernel_result_slice_4_valid => enable_passthrough_case_1_y_net_x4
  );
  result_muxer_5 : entity xil_defaultlib.mh_result_muxer_5 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    force_off => first_kernel_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_1_y_net_x3,
    kernel_result_slice_1_valid => enable_passthrough_case_1_y_net_x3,
    kernel_result_slice_2_valid => enable_passthrough_case_1_y_net_x3,
    kernel_result_slice_3_valid => enable_passthrough_case_1_y_net_x3,
    kernel_result_slice_4_valid => enable_passthrough_case_1_y_net_x3
  );
  result_muxer_6 : entity xil_defaultlib.mh_result_muxer_6 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    force_off => first_kernel_op_net,
    force_off_2 => last_kernel_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_1_y_net_x2,
    kernel_result_slice_1_valid => enable_passthrough_case_1_y_net_x2,
    kernel_result_slice_2_valid => enable_passthrough_case_1_y_net_x2,
    kernel_result_slice_3_valid => enable_passthrough_case_1_y_net_x2,
    kernel_result_slice_4_valid => enable_passthrough_case_0_y_net_x2
  );
  result_muxer_7 : entity xil_defaultlib.mh_result_muxer_7 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    force_off => first_kernel_op_net,
    force_off_2 => last_kernel_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_1_y_net_x1,
    kernel_result_slice_1_valid => enable_passthrough_case_1_y_net_x1,
    kernel_result_slice_2_valid => enable_passthrough_case_1_y_net_x1,
    kernel_result_slice_3_valid => enable_passthrough_case_0_y_net_x0,
    kernel_result_slice_4_valid => enable_passthrough_case_0_y_net_x0
  );
  result_muxer_8 : entity xil_defaultlib.mh_result_muxer_8 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    force_off => first_kernel_op_net,
    force_off_2 => last_kernel_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_1_y_net,
    kernel_result_slice_1_valid => enable_passthrough_case_1_y_net,
    kernel_result_slice_2_valid => enable_passthrough_case_0_y_net_x1,
    kernel_result_slice_3_valid => enable_passthrough_case_0_y_net_x1,
    kernel_result_slice_4_valid => enable_passthrough_case_0_y_net_x1
  );
  result_muxer_9 : entity xil_defaultlib.mh_result_muxer_9 
  port map (
    select_x0 => disable_q_net,
    valid => valid_data_delay_4_q_net,
    force_off => first_kernel_op_net,
    force_off_2 => last_kernel_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_slice_0_valid => enable_passthrough_case_1_y_net_x0,
    kernel_result_slice_1_valid => enable_passthrough_case_0_y_net,
    kernel_result_slice_2_valid => enable_passthrough_case_0_y_net,
    kernel_result_slice_3_valid => enable_passthrough_case_0_y_net,
    kernel_result_slice_4_valid => enable_passthrough_case_0_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_d5907f983e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  data_in : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 169,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i2",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    clr => '0',
    rst => valid_data_delay_6_q_net,
    en => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => data_in_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => relational1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  enable_disable_kernels : entity xil_defaultlib.sysgen_counter_4497493dc5 
  port map (
    clr => '0',
    rst => valid_data_delay_10_q_net,
    en => logical3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => enable_disable_kernels_op_net
  );
  enable_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_row_enable_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_delay2_q_net
  );
  disable : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_disable_kernels_op_net,
    clk => clk_net,
    ce => ce_net,
    q => disable_q_net
  );
  first_kernel : entity xil_defaultlib.sysgen_relational_f4134ca8cb 
  port map (
    clr => '0',
    a => constant_op_net,
    b => what_kernel_position_op_net,
    clk => clk_net,
    ce => ce_net,
    op => first_kernel_op_net
  );
  last_kernel_x0 : entity xil_defaultlib.sysgen_constant_13e8def457 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => last_kernel_op_net_x0
  );
  last_kernel : entity xil_defaultlib.sysgen_relational_5b9daf1b53 
  port map (
    clr => '0',
    a => what_kernel_position_op_net,
    b => last_kernel_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    op => last_kernel_op_net
  );
  last_out : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_out_q_net
  );
  last_row_enable_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => last_row_enable_delay_1_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => relational_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => data_valid_out_delay_q_net,
    d1 => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  logical2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => logical_y_net,
    d1 => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical2_y_net
  );
  logical3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => logical_y_net,
    d1 => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical3_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_665a4806e7 
  port map (
    clr => '0',
    a => data_in_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  relational1 : entity xil_defaultlib.sysgen_relational_6034f3e22a 
  port map (
    clr => '0',
    a => data_in_op_net,
    b => constant3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational1_op_net
  );
  valid_data_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_1_q_net
  );
  valid_data_delay_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_10_q_net
  );
  valid_data_delay_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_11_q_net
  );
  valid_data_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_2_q_net
  );
  valid_data_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_3_q_net
  );
  valid_data_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_4_q_net
  );
  valid_data_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => data_valid_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_5_q_net
  );
  valid_data_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_6_q_net
  );
  valid_data_delay_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => valid_data_delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_7_q_net
  );
  valid_data_delay_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => valid_data_delay_9_q_net
  );
  what_kernel_position : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 219,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i3",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 12
  )
  port map (
    clr => '0',
    rst => valid_data_delay_9_q_net,
    en => logical2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => what_kernel_position_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Organizer
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_organizer is
  port (
    in_pixel_0_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_weight_0_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    valid_data_in : in std_logic_vector( 1-1 downto 0 );
    reset_to_known_state : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    pixel_group_offset_0_1 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_1 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_1 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_1 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_1 : out std_logic_vector( 12-1 downto 0 );
    weights_1 : out std_logic_vector( 18-1 downto 0 );
    kernel_result_valid_bus_0_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_1_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_2_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_3_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_4_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_5_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_6_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_7_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_8_1 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_9_1 : out std_logic_vector( 1-1 downto 0 );
    pixel_group_offset_0_2 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_3 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_4 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_5 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_6 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_7 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_8 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_9 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_10 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_11 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_0_12 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_2 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_3 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_4 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_5 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_6 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_7 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_8 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_9 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_10 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_11 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_1_12 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_2 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_3 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_4 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_5 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_6 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_7 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_8 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_9 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_10 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_11 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_2_12 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_2 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_3 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_4 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_5 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_6 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_7 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_8 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_9 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_10 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_11 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_3_12 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_2 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_3 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_4 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_5 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_6 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_7 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_8 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_9 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_10 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_11 : out std_logic_vector( 12-1 downto 0 );
    pixel_group_offset_4_12 : out std_logic_vector( 12-1 downto 0 );
    weights_2 : out std_logic_vector( 18-1 downto 0 );
    weights_3 : out std_logic_vector( 18-1 downto 0 );
    weights_4 : out std_logic_vector( 18-1 downto 0 );
    weights_5 : out std_logic_vector( 18-1 downto 0 );
    weights_6 : out std_logic_vector( 18-1 downto 0 );
    weights_7 : out std_logic_vector( 18-1 downto 0 );
    weights_8 : out std_logic_vector( 18-1 downto 0 );
    weights_9 : out std_logic_vector( 18-1 downto 0 );
    weights_10 : out std_logic_vector( 18-1 downto 0 );
    weights_11 : out std_logic_vector( 18-1 downto 0 );
    weights_12 : out std_logic_vector( 18-1 downto 0 );
    weights_13 : out std_logic_vector( 18-1 downto 0 );
    weights_14 : out std_logic_vector( 18-1 downto 0 );
    weights_15 : out std_logic_vector( 18-1 downto 0 );
    weights_16 : out std_logic_vector( 18-1 downto 0 );
    weights_17 : out std_logic_vector( 18-1 downto 0 );
    weights_18 : out std_logic_vector( 18-1 downto 0 );
    weights_19 : out std_logic_vector( 18-1 downto 0 );
    weights_20 : out std_logic_vector( 18-1 downto 0 );
    weights_21 : out std_logic_vector( 18-1 downto 0 );
    weights_22 : out std_logic_vector( 18-1 downto 0 );
    weights_23 : out std_logic_vector( 18-1 downto 0 );
    weights_24 : out std_logic_vector( 18-1 downto 0 );
    weights_25 : out std_logic_vector( 18-1 downto 0 );
    weights_26 : out std_logic_vector( 18-1 downto 0 );
    weights_27 : out std_logic_vector( 18-1 downto 0 );
    weights_28 : out std_logic_vector( 18-1 downto 0 );
    weights_29 : out std_logic_vector( 18-1 downto 0 );
    weights_30 : out std_logic_vector( 18-1 downto 0 );
    weights_31 : out std_logic_vector( 18-1 downto 0 );
    weights_32 : out std_logic_vector( 18-1 downto 0 );
    weights_33 : out std_logic_vector( 18-1 downto 0 );
    weights_34 : out std_logic_vector( 18-1 downto 0 );
    weights_35 : out std_logic_vector( 18-1 downto 0 );
    weights_36 : out std_logic_vector( 18-1 downto 0 );
    weights_37 : out std_logic_vector( 18-1 downto 0 );
    weights_38 : out std_logic_vector( 18-1 downto 0 );
    weights_39 : out std_logic_vector( 18-1 downto 0 );
    weights_40 : out std_logic_vector( 18-1 downto 0 );
    weights_41 : out std_logic_vector( 18-1 downto 0 );
    weights_42 : out std_logic_vector( 18-1 downto 0 );
    weights_43 : out std_logic_vector( 18-1 downto 0 );
    weights_44 : out std_logic_vector( 18-1 downto 0 );
    weights_45 : out std_logic_vector( 18-1 downto 0 );
    weights_46 : out std_logic_vector( 18-1 downto 0 );
    weights_47 : out std_logic_vector( 18-1 downto 0 );
    weights_48 : out std_logic_vector( 18-1 downto 0 );
    weights_49 : out std_logic_vector( 18-1 downto 0 );
    weights_50 : out std_logic_vector( 18-1 downto 0 );
    weights_51 : out std_logic_vector( 18-1 downto 0 );
    weights_52 : out std_logic_vector( 18-1 downto 0 );
    weights_53 : out std_logic_vector( 18-1 downto 0 );
    weights_54 : out std_logic_vector( 18-1 downto 0 );
    weights_55 : out std_logic_vector( 18-1 downto 0 );
    weights_56 : out std_logic_vector( 18-1 downto 0 );
    weights_57 : out std_logic_vector( 18-1 downto 0 );
    weights_58 : out std_logic_vector( 18-1 downto 0 );
    weights_59 : out std_logic_vector( 18-1 downto 0 );
    weights_60 : out std_logic_vector( 18-1 downto 0 );
    weights_61 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_0_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_0_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_0_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_0_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_1_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_1_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_1_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_1_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_2_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_2_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_2_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_2_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_3_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_3_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_3_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_3_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_4_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_4_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_4_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_4_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_5_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_5_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_5_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_5_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_6_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_6_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_6_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_6_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_7_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_7_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_7_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_7_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_8_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_8_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_8_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_8_5 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_9_2 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_9_3 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_9_4 : out std_logic_vector( 1-1 downto 0 );
    kernel_result_valid_bus_9_5 : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_organizer;
architecture structural of mh_kernel_organizer is 
  signal delay_398_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_404_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_397_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_401_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_403_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_399_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_400_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_402_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_409_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_413_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_405_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_408_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_411_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_410_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_412_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_407_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_406_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_418_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_419_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_417_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_414_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_420_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_416_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_415_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_221_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_226_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_346_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_223_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_343_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_341_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_344_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_220_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_340_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_225_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_345_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_342_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_222_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_224_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_347_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_353_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_233_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_351_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_348_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_227_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_231_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_229_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_230_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_350_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_232_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_352_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_349_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_228_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_239_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_355_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_235_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_237_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_354_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_356_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_238_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_359_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_234_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_358_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_236_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_357_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_360_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_361_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_364_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_367_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_363_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_362_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_365_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_368_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_369_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_366_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_373_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_372_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_375_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_370_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_374_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_376_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_371_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_377_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_378_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_381_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_385_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_386_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_382_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_383_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_384_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_387_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_379_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_380_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_390_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_393_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_388_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_394_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_392_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_391_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_389_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_395_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_396_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_513_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_509_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_511_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_512_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_508_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_514_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_510_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_507_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_520_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_517_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_516_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_515_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_521_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_519_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_518_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_522_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_524_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_525_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_529_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_526_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_523_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_530_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_528_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_527_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_538_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_535_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_532_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_537_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_534_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_539_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_531_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_533_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_536_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_543_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_547_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_541_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_544_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_542_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_546_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_540_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_545_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_550_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_551_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_555_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_548_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_549_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_553_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_552_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_554_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_563_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_559_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_560_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_556_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_558_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_561_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_557_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_562_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_564_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_569_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_572_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_571_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_566_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_567_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_568_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_570_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_565_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_573_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_579_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_575_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_578_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_576_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_580_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_577_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_574_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_587_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_583_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_582_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_588_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_585_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_586_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_581_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_584_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_589_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_590_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_944_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_940_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_943_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_938_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_942_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_941_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_939_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_949_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_946_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_952_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_945_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_948_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_951_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_947_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_953_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_950_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_958_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_956_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_955_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_957_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_959_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_954_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_721_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_720_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_882_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_883_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_884_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_879_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_881_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_885_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_880_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_878_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_887_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_890_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_888_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_891_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_893_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_889_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_892_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_886_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_894_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_895_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_898_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_901_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_897_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_899_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_902_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_896_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_900_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_906_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_903_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_907_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_904_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_905_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_908_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_909_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_910_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_916_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_914_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_915_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_917_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_919_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_911_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_913_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_912_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_918_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_924_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_926_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_920_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_927_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_923_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_921_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_922_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_925_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_934_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_928_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_936_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_935_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_933_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_931_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_932_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_930_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_929_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_937_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_427_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_426_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_428_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_429_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_421_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_422_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_425_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_423_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_424_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_430_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_436_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_431_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_434_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_432_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_433_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_435_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_437_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_443_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_438_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_441_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_444_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_445_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_440_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_439_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_442_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_446_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_450_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_451_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_449_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_447_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_448_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_453_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_452_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_454_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_460_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_459_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_461_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_458_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_462_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_455_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_457_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_456_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_470_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_463_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_464_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_469_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_467_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_468_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_466_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_471_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_465_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_477_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_475_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_479_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_472_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_473_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_476_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_474_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_478_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_487_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_480_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_486_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_485_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_481_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_483_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_482_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_484_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_488_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_495_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_496_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_491_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_492_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_489_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_494_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_490_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_493_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_503_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_498_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_497_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_499_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_500_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_502_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_504_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_505_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_501_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_506_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_599_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_594_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_597_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_598_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_592_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_591_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_593_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_596_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_595_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_602_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_604_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_601_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_606_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_600_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_607_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_603_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_605_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_610_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_613_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_611_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_608_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_612_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_609_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_614_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_615_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_623_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_620_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_621_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_616_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_617_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_618_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_619_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_622_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_627_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_628_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_631_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_630_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_625_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_624_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_626_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_629_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_632_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_633_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_634_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_635_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_636_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_637_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_639_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_638_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_645_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_648_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_649_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_642_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_640_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_641_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_643_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_647_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_646_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_644_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_651_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_653_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_650_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_656_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_657_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_655_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_652_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_654_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_664_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_665_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_659_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_661_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_662_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_660_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_658_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_663_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_669_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_670_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_672_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_666_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_671_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_667_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_668_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_726_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_727_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_724_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_722_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_728_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_729_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_723_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_725_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_736_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_731_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_732_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_733_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_735_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_734_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_737_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_738_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_730_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_743_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_740_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_742_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_744_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_745_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_746_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_747_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_739_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_741_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_755_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_750_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_752_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_753_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_748_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_751_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_749_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_754_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_762_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_763_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_756_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_758_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_761_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_757_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_759_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_760_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_767_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_771_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_765_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_768_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_769_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_764_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_770_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_766_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_779_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_780_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_773_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_777_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_776_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_778_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_775_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_772_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_774_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_781_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_786_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_784_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_787_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_789_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_788_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_782_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_783_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_785_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_790_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_793_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_796_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_797_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_795_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_794_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_791_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_792_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_804_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_801_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_805_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_800_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_799_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_803_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_802_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_798_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_806_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_813_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_807_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_814_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_809_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_810_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_808_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_811_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_812_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_815_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_819_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_818_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_821_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_816_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_820_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_822_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_817_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_830_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_831_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_824_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_829_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_827_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_828_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_825_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_826_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_823_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_839_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_835_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_834_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_837_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_832_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_833_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_838_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_836_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_260_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_259_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_261_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_257_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_264_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_262_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_263_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_146_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_256_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_258_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_122_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_121_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_123_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_120_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_124_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal data_valid_out_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_130_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_127_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_126_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_128_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_131_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_129_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_132_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_125_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_133_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_141_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_137_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_134_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_140_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_135_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_139_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_142_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_138_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_136_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_144_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_244_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_243_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_143_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_245_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_240_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_246_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_241_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_242_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_250_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_252_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_251_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_249_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_145_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_248_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_253_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_254_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_247_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_255_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_873_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_876_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_874_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_877_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_875_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_870_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_871_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_869_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_872_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_677_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_679_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_675_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_674_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_680_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_676_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_678_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_673_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_686_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_688_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_681_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_689_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_683_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_684_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_682_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_685_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_687_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_695_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_698_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_696_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_692_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_691_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_690_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_693_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_694_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_697_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_705_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_699_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_703_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_700_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_706_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_701_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_702_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_704_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_711_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_709_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_710_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_712_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_708_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_707_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_713_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_714_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_842_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_715_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_717_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_718_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_840_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_841_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_719_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_716_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_847_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_850_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_845_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_843_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_846_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_848_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_849_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_844_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_851_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_857_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_859_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_853_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_855_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_852_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_854_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_856_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_858_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_860_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_862_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_867_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_865_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_863_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_864_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_861_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_866_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_868_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_269_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_268_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_267_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_147_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_149_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_266_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_150_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_270_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_265_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_148_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_151_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_271_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_159_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_275_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_276_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_279_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_152_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_156_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_153_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_154_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_157_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_273_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_277_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_155_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_272_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_274_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_278_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_158_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_164_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_280_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_281_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_282_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_283_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_165_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_285_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_162_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_284_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_160_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_161_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_163_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_166_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_286_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_294_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_289_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_290_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_287_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_169_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_171_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_170_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_292_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_172_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_173_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_168_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_167_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_293_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_291_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_174_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_288_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_175_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_298_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_295_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_178_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_299_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_297_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_181_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_300_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_177_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_179_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_180_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_301_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_176_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_296_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_189_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_183_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_304_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_303_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_187_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_307_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_188_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_308_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_302_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_306_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_185_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_182_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_305_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_186_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_184_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_309_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_195_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_315_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_313_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_316_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_312_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_194_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_191_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_311_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_314_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_310_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_196_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_192_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_193_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_190_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_203_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_323_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_199_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_197_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_317_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_319_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_318_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_198_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_200_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_320_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_321_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_202_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_322_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_201_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_326_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_329_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_204_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_205_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_327_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_210_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_207_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_325_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_206_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_324_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_330_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_209_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_208_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_328_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_216_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_337_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_214_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_334_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_217_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_335_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_215_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_213_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_332_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_218_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_338_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_336_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_211_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_212_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_333_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_331_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_339_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_219_q_net : std_logic_vector( 12-1 downto 0 );
begin
  pixel_group_offset_0_1 <= delay_0_q_net;
  pixel_group_offset_1_1 <= delay_22_q_net;
  pixel_group_offset_2_1 <= delay_48_q_net;
  pixel_group_offset_3_1 <= delay_72_q_net;
  pixel_group_offset_4_1 <= delay_96_q_net;
  weights_1 <= delay_1_q_net;
  kernel_result_valid_bus_0_1 <= enable_passthrough_case_0_y_net;
  kernel_result_valid_bus_1_1 <= enable_passthrough_case_0_y_net_x0;
  kernel_result_valid_bus_2_1 <= enable_passthrough_case_0_y_net_x1;
  kernel_result_valid_bus_3_1 <= enable_passthrough_case_0_y_net_x2;
  kernel_result_valid_bus_4_1 <= enable_passthrough_case_0_y_net_x3;
  kernel_result_valid_bus_5_1 <= enable_passthrough_case_1_y_net_x3;
  kernel_result_valid_bus_6_1 <= enable_passthrough_case_1_y_net_x4;
  kernel_result_valid_bus_7_1 <= enable_passthrough_case_1_y_net_x5;
  kernel_result_valid_bus_8_1 <= enable_passthrough_case_1_y_net_x6;
  kernel_result_valid_bus_9_1 <= enable_passthrough_case_1_y_net_x7;
  pixel_group_offset_0_2 <= delay_2_q_net;
  pixel_group_offset_0_3 <= delay_4_q_net;
  pixel_group_offset_0_4 <= delay_6_q_net;
  pixel_group_offset_0_5 <= delay_8_q_net;
  pixel_group_offset_0_6 <= delay_10_q_net;
  pixel_group_offset_0_7 <= delay_12_q_net;
  pixel_group_offset_0_8 <= delay_14_q_net;
  pixel_group_offset_0_9 <= delay_23_q_net;
  pixel_group_offset_0_10 <= delay_16_q_net;
  pixel_group_offset_0_11 <= delay_18_q_net;
  pixel_group_offset_0_12 <= delay_20_q_net;
  pixel_group_offset_1_2 <= delay_36_q_net;
  pixel_group_offset_1_3 <= delay_42_q_net;
  pixel_group_offset_1_4 <= delay_44_q_net;
  pixel_group_offset_1_5 <= delay_46_q_net;
  pixel_group_offset_1_6 <= delay_26_q_net;
  pixel_group_offset_1_7 <= delay_28_q_net;
  pixel_group_offset_1_8 <= delay_30_q_net;
  pixel_group_offset_1_9 <= delay_39_q_net;
  pixel_group_offset_1_10 <= delay_32_q_net;
  pixel_group_offset_1_11 <= delay_34_q_net;
  pixel_group_offset_1_12 <= delay_37_q_net;
  pixel_group_offset_2_2 <= delay_60_q_net;
  pixel_group_offset_2_3 <= delay_66_q_net;
  pixel_group_offset_2_4 <= delay_68_q_net;
  pixel_group_offset_2_5 <= delay_70_q_net;
  pixel_group_offset_2_6 <= delay_50_q_net;
  pixel_group_offset_2_7 <= delay_52_q_net;
  pixel_group_offset_2_8 <= delay_54_q_net;
  pixel_group_offset_2_9 <= delay_63_q_net;
  pixel_group_offset_2_10 <= delay_56_q_net;
  pixel_group_offset_2_11 <= delay_58_q_net;
  pixel_group_offset_2_12 <= delay_61_q_net;
  pixel_group_offset_3_2 <= delay_84_q_net;
  pixel_group_offset_3_3 <= delay_90_q_net;
  pixel_group_offset_3_4 <= delay_92_q_net;
  pixel_group_offset_3_5 <= delay_94_q_net;
  pixel_group_offset_3_6 <= delay_74_q_net;
  pixel_group_offset_3_7 <= delay_76_q_net;
  pixel_group_offset_3_8 <= delay_78_q_net;
  pixel_group_offset_3_9 <= delay_87_q_net;
  pixel_group_offset_3_10 <= delay_80_q_net;
  pixel_group_offset_3_11 <= delay_82_q_net;
  pixel_group_offset_3_12 <= delay_85_q_net;
  pixel_group_offset_4_2 <= delay_108_q_net;
  pixel_group_offset_4_3 <= delay_114_q_net;
  pixel_group_offset_4_4 <= delay_116_q_net;
  pixel_group_offset_4_5 <= delay_118_q_net;
  pixel_group_offset_4_6 <= delay_98_q_net;
  pixel_group_offset_4_7 <= delay_100_q_net;
  pixel_group_offset_4_8 <= delay_102_q_net;
  pixel_group_offset_4_9 <= delay_111_q_net;
  pixel_group_offset_4_10 <= delay_104_q_net;
  pixel_group_offset_4_11 <= delay_106_q_net;
  pixel_group_offset_4_12 <= delay_109_q_net;
  weights_2 <= delay_3_q_net;
  weights_3 <= delay_5_q_net;
  weights_4 <= delay_7_q_net;
  weights_5 <= delay_9_q_net;
  weights_6 <= delay_11_q_net;
  weights_7 <= delay_13_q_net;
  weights_8 <= delay_15_q_net;
  weights_9 <= delay_24_q_net;
  weights_10 <= delay_17_q_net;
  weights_11 <= delay_19_q_net;
  weights_12 <= delay_21_q_net;
  weights_13 <= delay_25_q_net;
  weights_14 <= delay_41_q_net;
  weights_15 <= delay_43_q_net;
  weights_16 <= delay_45_q_net;
  weights_17 <= delay_47_q_net;
  weights_18 <= delay_27_q_net;
  weights_19 <= delay_29_q_net;
  weights_20 <= delay_31_q_net;
  weights_21 <= delay_40_q_net;
  weights_22 <= delay_33_q_net;
  weights_23 <= delay_35_q_net;
  weights_24 <= delay_38_q_net;
  weights_25 <= delay_49_q_net;
  weights_26 <= delay_65_q_net;
  weights_27 <= delay_67_q_net;
  weights_28 <= delay_69_q_net;
  weights_29 <= delay_71_q_net;
  weights_30 <= delay_51_q_net;
  weights_31 <= delay_53_q_net;
  weights_32 <= delay_55_q_net;
  weights_33 <= delay_64_q_net;
  weights_34 <= delay_57_q_net;
  weights_35 <= delay_59_q_net;
  weights_36 <= delay_62_q_net;
  weights_37 <= delay_73_q_net;
  weights_38 <= delay_89_q_net;
  weights_39 <= delay_91_q_net;
  weights_40 <= delay_93_q_net;
  weights_41 <= delay_95_q_net;
  weights_42 <= delay_75_q_net;
  weights_43 <= delay_77_q_net;
  weights_44 <= delay_79_q_net;
  weights_45 <= delay_88_q_net;
  weights_46 <= delay_81_q_net;
  weights_47 <= delay_83_q_net;
  weights_48 <= delay_86_q_net;
  weights_49 <= delay_97_q_net;
  weights_50 <= delay_113_q_net;
  weights_51 <= delay_115_q_net;
  weights_52 <= delay_117_q_net;
  weights_53 <= delay_119_q_net;
  weights_54 <= delay_99_q_net;
  weights_55 <= delay_101_q_net;
  weights_56 <= delay_103_q_net;
  weights_57 <= delay_112_q_net;
  weights_58 <= delay_105_q_net;
  weights_59 <= delay_107_q_net;
  weights_60 <= delay_110_q_net;
  weights_61 <= last_out_q_net;
  kernel_result_valid_bus_0_2 <= enable_passthrough_case_0_y_net;
  kernel_result_valid_bus_0_3 <= enable_passthrough_case_0_y_net;
  kernel_result_valid_bus_0_4 <= enable_passthrough_case_0_y_net;
  kernel_result_valid_bus_0_5 <= enable_passthrough_case_0_y_net;
  kernel_result_valid_bus_1_2 <= enable_passthrough_case_0_y_net_x0;
  kernel_result_valid_bus_1_3 <= enable_passthrough_case_0_y_net_x0;
  kernel_result_valid_bus_1_4 <= enable_passthrough_case_0_y_net_x0;
  kernel_result_valid_bus_1_5 <= enable_passthrough_case_1_y_net;
  kernel_result_valid_bus_2_2 <= enable_passthrough_case_0_y_net_x1;
  kernel_result_valid_bus_2_3 <= enable_passthrough_case_0_y_net_x1;
  kernel_result_valid_bus_2_4 <= enable_passthrough_case_1_y_net_x0;
  kernel_result_valid_bus_2_5 <= enable_passthrough_case_1_y_net_x0;
  kernel_result_valid_bus_3_2 <= enable_passthrough_case_0_y_net_x2;
  kernel_result_valid_bus_3_3 <= enable_passthrough_case_1_y_net_x1;
  kernel_result_valid_bus_3_4 <= enable_passthrough_case_1_y_net_x1;
  kernel_result_valid_bus_3_5 <= enable_passthrough_case_1_y_net_x1;
  kernel_result_valid_bus_4_2 <= enable_passthrough_case_1_y_net_x2;
  kernel_result_valid_bus_4_3 <= enable_passthrough_case_1_y_net_x2;
  kernel_result_valid_bus_4_4 <= enable_passthrough_case_1_y_net_x2;
  kernel_result_valid_bus_4_5 <= enable_passthrough_case_1_y_net_x2;
  kernel_result_valid_bus_5_2 <= enable_passthrough_case_1_y_net_x3;
  kernel_result_valid_bus_5_3 <= enable_passthrough_case_1_y_net_x3;
  kernel_result_valid_bus_5_4 <= enable_passthrough_case_1_y_net_x3;
  kernel_result_valid_bus_5_5 <= enable_passthrough_case_1_y_net_x3;
  kernel_result_valid_bus_6_2 <= enable_passthrough_case_1_y_net_x4;
  kernel_result_valid_bus_6_3 <= enable_passthrough_case_1_y_net_x4;
  kernel_result_valid_bus_6_4 <= enable_passthrough_case_1_y_net_x4;
  kernel_result_valid_bus_6_5 <= enable_passthrough_case_0_y_net_x4;
  kernel_result_valid_bus_7_2 <= enable_passthrough_case_1_y_net_x5;
  kernel_result_valid_bus_7_3 <= enable_passthrough_case_1_y_net_x5;
  kernel_result_valid_bus_7_4 <= enable_passthrough_case_0_y_net_x5;
  kernel_result_valid_bus_7_5 <= enable_passthrough_case_0_y_net_x5;
  kernel_result_valid_bus_8_2 <= enable_passthrough_case_1_y_net_x6;
  kernel_result_valid_bus_8_3 <= enable_passthrough_case_0_y_net_x6;
  kernel_result_valid_bus_8_4 <= enable_passthrough_case_0_y_net_x6;
  kernel_result_valid_bus_8_5 <= enable_passthrough_case_0_y_net_x6;
  kernel_result_valid_bus_9_2 <= enable_passthrough_case_0_y_net_x7;
  kernel_result_valid_bus_9_3 <= enable_passthrough_case_0_y_net_x7;
  kernel_result_valid_bus_9_4 <= enable_passthrough_case_0_y_net_x7;
  kernel_result_valid_bus_9_5 <= enable_passthrough_case_0_y_net_x7;
  x12_bit_bin_value_0_q_net_x8 <= in_pixel_0_at_offset_0;
  x12_bit_bin_value_1_q_net_x8 <= in_pixel_1_at_offset_0;
  x12_bit_bin_value_2_q_net_x8 <= in_pixel_2_at_offset_0;
  x12_bit_bin_value_3_q_net_x8 <= in_pixel_3_at_offset_0;
  x12_bit_bin_value_4_q_net_x8 <= in_pixel_4_at_offset_0;
  x12_bit_bin_value_5_q_net_x8 <= in_pixel_5_at_offset_0;
  x12_bit_bin_value_6_q_net_x8 <= in_pixel_6_at_offset_0;
  x12_bit_bin_value_7_q_net_x8 <= in_pixel_7_at_offset_0;
  x12_bit_bin_value_8_q_net_x8 <= in_pixel_8_at_offset_0;
  x12_bit_bin_value_9_q_net_x8 <= in_pixel_9_at_offset_0;
  x12_bit_bin_value_10_q_net_x8 <= in_pixel_10_at_offset_0;
  x12_bit_bin_value_11_q_net_x8 <= in_pixel_11_at_offset_0;
  x12_bit_bin_value_0_q_net_x7 <= in_pixel_0_at_offset_1;
  x12_bit_bin_value_1_q_net_x7 <= in_pixel_1_at_offset_1;
  x12_bit_bin_value_2_q_net_x7 <= in_pixel_2_at_offset_1;
  x12_bit_bin_value_3_q_net_x7 <= in_pixel_3_at_offset_1;
  x12_bit_bin_value_4_q_net_x7 <= in_pixel_4_at_offset_1;
  x12_bit_bin_value_5_q_net_x7 <= in_pixel_5_at_offset_1;
  x12_bit_bin_value_6_q_net_x7 <= in_pixel_6_at_offset_1;
  x12_bit_bin_value_7_q_net_x7 <= in_pixel_7_at_offset_1;
  x12_bit_bin_value_8_q_net_x7 <= in_pixel_8_at_offset_1;
  x12_bit_bin_value_9_q_net_x7 <= in_pixel_9_at_offset_1;
  x12_bit_bin_value_10_q_net_x7 <= in_pixel_10_at_offset_1;
  x12_bit_bin_value_11_q_net_x7 <= in_pixel_11_at_offset_1;
  x12_bit_bin_value_0_q_net_x6 <= in_pixel_0_at_offset_2;
  x12_bit_bin_value_1_q_net_x6 <= in_pixel_1_at_offset_2;
  x12_bit_bin_value_2_q_net_x6 <= in_pixel_2_at_offset_2;
  x12_bit_bin_value_3_q_net_x6 <= in_pixel_3_at_offset_2;
  x12_bit_bin_value_4_q_net_x6 <= in_pixel_4_at_offset_2;
  x12_bit_bin_value_5_q_net_x6 <= in_pixel_5_at_offset_2;
  x12_bit_bin_value_6_q_net_x6 <= in_pixel_6_at_offset_2;
  x12_bit_bin_value_7_q_net_x6 <= in_pixel_7_at_offset_2;
  x12_bit_bin_value_8_q_net_x6 <= in_pixel_8_at_offset_2;
  x12_bit_bin_value_9_q_net_x6 <= in_pixel_9_at_offset_2;
  x12_bit_bin_value_10_q_net_x6 <= in_pixel_10_at_offset_2;
  x12_bit_bin_value_11_q_net_x6 <= in_pixel_11_at_offset_2;
  x12_bit_bin_value_0_q_net_x5 <= in_pixel_0_at_offset_3;
  x12_bit_bin_value_1_q_net_x5 <= in_pixel_1_at_offset_3;
  x12_bit_bin_value_2_q_net_x5 <= in_pixel_2_at_offset_3;
  x12_bit_bin_value_3_q_net_x5 <= in_pixel_3_at_offset_3;
  x12_bit_bin_value_4_q_net_x5 <= in_pixel_4_at_offset_3;
  x12_bit_bin_value_5_q_net_x5 <= in_pixel_5_at_offset_3;
  x12_bit_bin_value_6_q_net_x5 <= in_pixel_6_at_offset_3;
  x12_bit_bin_value_7_q_net_x5 <= in_pixel_7_at_offset_3;
  x12_bit_bin_value_8_q_net_x5 <= in_pixel_8_at_offset_3;
  x12_bit_bin_value_9_q_net_x5 <= in_pixel_9_at_offset_3;
  x12_bit_bin_value_10_q_net_x5 <= in_pixel_10_at_offset_3;
  x12_bit_bin_value_11_q_net_x5 <= in_pixel_11_at_offset_3;
  x12_bit_bin_value_0_q_net_x4 <= in_pixel_0_at_offset_4;
  x12_bit_bin_value_1_q_net_x4 <= in_pixel_1_at_offset_4;
  x12_bit_bin_value_2_q_net_x4 <= in_pixel_2_at_offset_4;
  x12_bit_bin_value_3_q_net_x4 <= in_pixel_3_at_offset_4;
  x12_bit_bin_value_4_q_net_x4 <= in_pixel_4_at_offset_4;
  x12_bit_bin_value_5_q_net_x4 <= in_pixel_5_at_offset_4;
  x12_bit_bin_value_6_q_net_x4 <= in_pixel_6_at_offset_4;
  x12_bit_bin_value_7_q_net_x4 <= in_pixel_7_at_offset_4;
  x12_bit_bin_value_8_q_net_x4 <= in_pixel_8_at_offset_4;
  x12_bit_bin_value_9_q_net_x4 <= in_pixel_9_at_offset_4;
  x12_bit_bin_value_10_q_net_x4 <= in_pixel_10_at_offset_4;
  x12_bit_bin_value_11_q_net_x4 <= in_pixel_11_at_offset_4;
  x12_bit_bin_value_0_q_net_x3 <= in_weight_0_at_offset_0;
  x12_bit_bin_value_1_q_net_x3 <= in_weight_1_at_offset_0;
  x12_bit_bin_value_2_q_net_x3 <= in_weight_2_at_offset_0;
  x12_bit_bin_value_3_q_net_x3 <= in_weight_3_at_offset_0;
  x12_bit_bin_value_4_q_net_x3 <= in_weight_4_at_offset_0;
  x12_bit_bin_value_5_q_net_x3 <= in_weight_5_at_offset_0;
  x12_bit_bin_value_6_q_net_x3 <= in_weight_6_at_offset_0;
  x12_bit_bin_value_7_q_net_x3 <= in_weight_7_at_offset_0;
  x12_bit_bin_value_8_q_net_x3 <= in_weight_8_at_offset_0;
  x12_bit_bin_value_9_q_net_x3 <= in_weight_9_at_offset_0;
  x12_bit_bin_value_10_q_net_x3 <= in_weight_10_at_offset_0;
  x12_bit_bin_value_11_q_net_x3 <= in_weight_11_at_offset_0;
  x12_bit_bin_value_0_q_net_x2 <= in_weight_0_at_offset_1;
  x12_bit_bin_value_1_q_net_x2 <= in_weight_1_at_offset_1;
  x12_bit_bin_value_2_q_net_x2 <= in_weight_2_at_offset_1;
  x12_bit_bin_value_3_q_net_x2 <= in_weight_3_at_offset_1;
  x12_bit_bin_value_4_q_net_x2 <= in_weight_4_at_offset_1;
  x12_bit_bin_value_5_q_net_x2 <= in_weight_5_at_offset_1;
  x12_bit_bin_value_6_q_net_x2 <= in_weight_6_at_offset_1;
  x12_bit_bin_value_7_q_net_x2 <= in_weight_7_at_offset_1;
  x12_bit_bin_value_8_q_net_x2 <= in_weight_8_at_offset_1;
  x12_bit_bin_value_9_q_net_x2 <= in_weight_9_at_offset_1;
  x12_bit_bin_value_10_q_net_x2 <= in_weight_10_at_offset_1;
  x12_bit_bin_value_11_q_net_x2 <= in_weight_11_at_offset_1;
  x12_bit_bin_value_0_q_net_x1 <= in_weight_0_at_offset_2;
  x12_bit_bin_value_1_q_net_x1 <= in_weight_1_at_offset_2;
  x12_bit_bin_value_2_q_net_x1 <= in_weight_2_at_offset_2;
  x12_bit_bin_value_3_q_net_x1 <= in_weight_3_at_offset_2;
  x12_bit_bin_value_4_q_net_x1 <= in_weight_4_at_offset_2;
  x12_bit_bin_value_5_q_net_x1 <= in_weight_5_at_offset_2;
  x12_bit_bin_value_6_q_net_x1 <= in_weight_6_at_offset_2;
  x12_bit_bin_value_7_q_net_x1 <= in_weight_7_at_offset_2;
  x12_bit_bin_value_8_q_net_x1 <= in_weight_8_at_offset_2;
  x12_bit_bin_value_9_q_net_x1 <= in_weight_9_at_offset_2;
  x12_bit_bin_value_10_q_net_x1 <= in_weight_10_at_offset_2;
  x12_bit_bin_value_11_q_net_x1 <= in_weight_11_at_offset_2;
  x12_bit_bin_value_0_q_net_x0 <= in_weight_0_at_offset_3;
  x12_bit_bin_value_1_q_net_x0 <= in_weight_1_at_offset_3;
  x12_bit_bin_value_2_q_net_x0 <= in_weight_2_at_offset_3;
  x12_bit_bin_value_3_q_net_x0 <= in_weight_3_at_offset_3;
  x12_bit_bin_value_4_q_net_x0 <= in_weight_4_at_offset_3;
  x12_bit_bin_value_5_q_net_x0 <= in_weight_5_at_offset_3;
  x12_bit_bin_value_6_q_net_x0 <= in_weight_6_at_offset_3;
  x12_bit_bin_value_7_q_net_x0 <= in_weight_7_at_offset_3;
  x12_bit_bin_value_8_q_net_x0 <= in_weight_8_at_offset_3;
  x12_bit_bin_value_9_q_net_x0 <= in_weight_9_at_offset_3;
  x12_bit_bin_value_10_q_net_x0 <= in_weight_10_at_offset_3;
  x12_bit_bin_value_11_q_net_x0 <= in_weight_11_at_offset_3;
  x12_bit_bin_value_0_q_net <= in_weight_0_at_offset_4;
  x12_bit_bin_value_1_q_net <= in_weight_1_at_offset_4;
  x12_bit_bin_value_2_q_net <= in_weight_2_at_offset_4;
  x12_bit_bin_value_3_q_net <= in_weight_3_at_offset_4;
  x12_bit_bin_value_4_q_net <= in_weight_4_at_offset_4;
  x12_bit_bin_value_5_q_net <= in_weight_5_at_offset_4;
  x12_bit_bin_value_6_q_net <= in_weight_6_at_offset_4;
  x12_bit_bin_value_7_q_net <= in_weight_7_at_offset_4;
  x12_bit_bin_value_8_q_net <= in_weight_8_at_offset_4;
  x12_bit_bin_value_9_q_net <= in_weight_9_at_offset_4;
  x12_bit_bin_value_10_q_net <= in_weight_10_at_offset_4;
  x12_bit_bin_value_11_q_net <= in_weight_11_at_offset_4;
  data_valid_out_delay_q_net <= valid_data_in;
  switch_to_zero_y_net <= reset_to_known_state;
  clk_net <= clk_1;
  ce_net <= ce_1;
  determine_calculations_delay_1 : entity xil_defaultlib.mh_determine_calculations_delay_1 
  port map (
    valid_data_in => data_valid_out_delay_q_net,
    hard_reset => switch_to_zero_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_valid_out_0_kernel_result_0 => enable_passthrough_case_0_y_net,
    slice_valid_out_1_kernel_result_0 => enable_passthrough_case_0_y_net,
    slice_valid_out_2_kernel_result_0 => enable_passthrough_case_0_y_net,
    slice_valid_out_3_kernel_result_0 => enable_passthrough_case_0_y_net,
    slice_valid_out_4_kernel_result_0 => enable_passthrough_case_0_y_net,
    slice_valid_out_0_kernel_result_1 => enable_passthrough_case_0_y_net_x0,
    slice_valid_out_1_kernel_result_1 => enable_passthrough_case_0_y_net_x0,
    slice_valid_out_2_kernel_result_1 => enable_passthrough_case_0_y_net_x0,
    slice_valid_out_3_kernel_result_1 => enable_passthrough_case_0_y_net_x0,
    slice_valid_out_4_kernel_result_1 => enable_passthrough_case_1_y_net,
    slice_valid_out_0_kernel_result_2 => enable_passthrough_case_0_y_net_x1,
    slice_valid_out_1_kernel_result_2 => enable_passthrough_case_0_y_net_x1,
    slice_valid_out_2_kernel_result_2 => enable_passthrough_case_0_y_net_x1,
    slice_valid_out_3_kernel_result_2 => enable_passthrough_case_1_y_net_x0,
    slice_valid_out_4_kernel_result_2 => enable_passthrough_case_1_y_net_x0,
    slice_valid_out_0_kernel_result_3 => enable_passthrough_case_0_y_net_x2,
    slice_valid_out_1_kernel_result_3 => enable_passthrough_case_0_y_net_x2,
    slice_valid_out_2_kernel_result_3 => enable_passthrough_case_1_y_net_x1,
    slice_valid_out_3_kernel_result_3 => enable_passthrough_case_1_y_net_x1,
    slice_valid_out_4_kernel_result_3 => enable_passthrough_case_1_y_net_x1,
    slice_valid_out_0_kernel_result_4 => enable_passthrough_case_0_y_net_x3,
    slice_valid_out_1_kernel_result_4 => enable_passthrough_case_1_y_net_x2,
    slice_valid_out_2_kernel_result_4 => enable_passthrough_case_1_y_net_x2,
    slice_valid_out_3_kernel_result_4 => enable_passthrough_case_1_y_net_x2,
    slice_valid_out_4_kernel_result_4 => enable_passthrough_case_1_y_net_x2,
    slice_valid_out_0_kernel_result_5 => enable_passthrough_case_1_y_net_x3,
    slice_valid_out_1_kernel_result_5 => enable_passthrough_case_1_y_net_x3,
    slice_valid_out_2_kernel_result_5 => enable_passthrough_case_1_y_net_x3,
    slice_valid_out_3_kernel_result_5 => enable_passthrough_case_1_y_net_x3,
    slice_valid_out_4_kernel_result_5 => enable_passthrough_case_1_y_net_x3,
    slice_valid_out_0_kernel_result_6 => enable_passthrough_case_1_y_net_x4,
    slice_valid_out_1_kernel_result_6 => enable_passthrough_case_1_y_net_x4,
    slice_valid_out_2_kernel_result_6 => enable_passthrough_case_1_y_net_x4,
    slice_valid_out_3_kernel_result_6 => enable_passthrough_case_1_y_net_x4,
    slice_valid_out_4_kernel_result_6 => enable_passthrough_case_0_y_net_x4,
    slice_valid_out_0_kernel_result_7 => enable_passthrough_case_1_y_net_x5,
    slice_valid_out_1_kernel_result_7 => enable_passthrough_case_1_y_net_x5,
    slice_valid_out_2_kernel_result_7 => enable_passthrough_case_1_y_net_x5,
    slice_valid_out_3_kernel_result_7 => enable_passthrough_case_0_y_net_x5,
    slice_valid_out_4_kernel_result_7 => enable_passthrough_case_0_y_net_x5,
    slice_valid_out_0_kernel_result_8 => enable_passthrough_case_1_y_net_x6,
    slice_valid_out_1_kernel_result_8 => enable_passthrough_case_1_y_net_x6,
    slice_valid_out_2_kernel_result_8 => enable_passthrough_case_0_y_net_x6,
    slice_valid_out_3_kernel_result_8 => enable_passthrough_case_0_y_net_x6,
    slice_valid_out_4_kernel_result_8 => enable_passthrough_case_0_y_net_x6,
    slice_valid_out_0_kernel_result_9 => enable_passthrough_case_1_y_net_x7,
    slice_valid_out_1_kernel_result_9 => enable_passthrough_case_0_y_net_x7,
    slice_valid_out_2_kernel_result_9 => enable_passthrough_case_0_y_net_x7,
    slice_valid_out_3_kernel_result_9 => enable_passthrough_case_0_y_net_x7,
    slice_valid_out_4_kernel_result_9 => enable_passthrough_case_0_y_net_x7,
    slice_valid_out_0_kernel_result_10 => last_out_q_net
  );
  delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_120_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_0_q_net
  );
  delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_121_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_1_q_net
  );
  delay_10 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_122_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_10_q_net
  );
  delay_100 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_123_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_100_q_net
  );
  delay_101 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_124_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_101_q_net
  );
  delay_102 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_125_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_102_q_net
  );
  delay_103 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_126_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_103_q_net
  );
  delay_104 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_127_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_104_q_net
  );
  delay_105 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_128_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_105_q_net
  );
  delay_106 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_129_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_106_q_net
  );
  delay_107 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_130_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_107_q_net
  );
  delay_108 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_131_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_108_q_net
  );
  delay_109 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_132_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_109_q_net
  );
  delay_11 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_133_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_11_q_net
  );
  delay_110 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_134_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_110_q_net
  );
  delay_111 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_135_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_111_q_net
  );
  delay_112 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_136_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_112_q_net
  );
  delay_113 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_137_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_113_q_net
  );
  delay_114 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_138_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_114_q_net
  );
  delay_115 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_139_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_115_q_net
  );
  delay_116 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_140_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_116_q_net
  );
  delay_117 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_141_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_117_q_net
  );
  delay_118 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_142_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_118_q_net
  );
  delay_119 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_143_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_119_q_net
  );
  delay_12 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_144_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_12_q_net
  );
  delay_120 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_240_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_120_q_net
  );
  delay_121 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_241_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_121_q_net
  );
  delay_122 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_242_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_122_q_net
  );
  delay_123 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_243_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_123_q_net
  );
  delay_124 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_244_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_124_q_net
  );
  delay_125 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_245_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_125_q_net
  );
  delay_126 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_246_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_126_q_net
  );
  delay_127 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_247_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_127_q_net
  );
  delay_128 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_248_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_128_q_net
  );
  delay_129 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_249_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_129_q_net
  );
  delay_13 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_145_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_13_q_net
  );
  delay_130 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_250_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_130_q_net
  );
  delay_131 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_251_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_131_q_net
  );
  delay_132 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_252_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_132_q_net
  );
  delay_133 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_253_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_133_q_net
  );
  delay_134 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_254_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_134_q_net
  );
  delay_135 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_255_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_135_q_net
  );
  delay_136 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_256_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_136_q_net
  );
  delay_137 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_257_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_137_q_net
  );
  delay_138 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_258_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_138_q_net
  );
  delay_139 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_259_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_139_q_net
  );
  delay_14 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_146_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_14_q_net
  );
  delay_140 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_260_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_140_q_net
  );
  delay_141 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_261_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_141_q_net
  );
  delay_142 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_262_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_142_q_net
  );
  delay_143 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_263_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_143_q_net
  );
  delay_144 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_264_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_144_q_net
  );
  delay_145 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_265_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_145_q_net
  );
  delay_146 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_266_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_146_q_net
  );
  delay_147 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_267_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_147_q_net
  );
  delay_148 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_268_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_148_q_net
  );
  delay_149 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_269_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_149_q_net
  );
  delay_15 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_147_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_15_q_net
  );
  delay_150 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_270_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_150_q_net
  );
  delay_151 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_271_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_151_q_net
  );
  delay_152 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_272_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_152_q_net
  );
  delay_153 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_273_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_153_q_net
  );
  delay_154 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_274_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_154_q_net
  );
  delay_155 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_275_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_155_q_net
  );
  delay_156 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_276_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_156_q_net
  );
  delay_157 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_277_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_157_q_net
  );
  delay_158 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_278_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_158_q_net
  );
  delay_159 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_279_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_159_q_net
  );
  delay_16 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_148_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_16_q_net
  );
  delay_160 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_280_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_160_q_net
  );
  delay_161 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_281_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_161_q_net
  );
  delay_162 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_282_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_162_q_net
  );
  delay_163 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_283_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_163_q_net
  );
  delay_164 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_284_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_164_q_net
  );
  delay_165 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_285_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_165_q_net
  );
  delay_166 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_286_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_166_q_net
  );
  delay_167 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_287_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_167_q_net
  );
  delay_168 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_288_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_168_q_net
  );
  delay_169 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_289_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_169_q_net
  );
  delay_17 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_149_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_17_q_net
  );
  delay_170 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_290_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_170_q_net
  );
  delay_171 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_291_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_171_q_net
  );
  delay_172 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_292_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_172_q_net
  );
  delay_173 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_293_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_173_q_net
  );
  delay_174 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_294_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_174_q_net
  );
  delay_175 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_295_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_175_q_net
  );
  delay_176 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_296_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_176_q_net
  );
  delay_177 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_297_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_177_q_net
  );
  delay_178 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_298_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_178_q_net
  );
  delay_179 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_299_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_179_q_net
  );
  delay_18 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_150_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_18_q_net
  );
  delay_180 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_300_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_180_q_net
  );
  delay_181 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_301_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_181_q_net
  );
  delay_182 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_302_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_182_q_net
  );
  delay_183 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_303_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_183_q_net
  );
  delay_184 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_304_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_184_q_net
  );
  delay_185 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_305_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_185_q_net
  );
  delay_186 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_306_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_186_q_net
  );
  delay_187 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_307_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_187_q_net
  );
  delay_188 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_308_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_188_q_net
  );
  delay_189 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_309_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_189_q_net
  );
  delay_19 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_151_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_19_q_net
  );
  delay_190 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_310_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_190_q_net
  );
  delay_191 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_311_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_191_q_net
  );
  delay_192 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_312_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_192_q_net
  );
  delay_193 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_313_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_193_q_net
  );
  delay_194 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_314_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_194_q_net
  );
  delay_195 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_315_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_195_q_net
  );
  delay_196 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_316_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_196_q_net
  );
  delay_197 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_317_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_197_q_net
  );
  delay_198 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_318_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_198_q_net
  );
  delay_199 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_319_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_199_q_net
  );
  delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_152_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_2_q_net
  );
  delay_20 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_153_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_20_q_net
  );
  delay_200 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_320_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_200_q_net
  );
  delay_201 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_321_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_201_q_net
  );
  delay_202 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_322_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_202_q_net
  );
  delay_203 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_323_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_203_q_net
  );
  delay_204 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_324_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_204_q_net
  );
  delay_205 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_325_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_205_q_net
  );
  delay_206 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_326_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_206_q_net
  );
  delay_207 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_327_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_207_q_net
  );
  delay_208 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_328_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_208_q_net
  );
  delay_209 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_329_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_209_q_net
  );
  delay_21 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_154_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_21_q_net
  );
  delay_210 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_330_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_210_q_net
  );
  delay_211 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_331_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_211_q_net
  );
  delay_212 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_332_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_212_q_net
  );
  delay_213 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_333_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_213_q_net
  );
  delay_214 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_334_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_214_q_net
  );
  delay_215 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_335_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_215_q_net
  );
  delay_216 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_336_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_216_q_net
  );
  delay_217 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_337_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_217_q_net
  );
  delay_218 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_338_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_218_q_net
  );
  delay_219 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_339_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_219_q_net
  );
  delay_22 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_155_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_22_q_net
  );
  delay_220 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_340_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_220_q_net
  );
  delay_221 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_341_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_221_q_net
  );
  delay_222 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_342_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_222_q_net
  );
  delay_223 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_343_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_223_q_net
  );
  delay_224 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_344_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_224_q_net
  );
  delay_225 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_345_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_225_q_net
  );
  delay_226 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_346_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_226_q_net
  );
  delay_227 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_347_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_227_q_net
  );
  delay_228 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_348_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_228_q_net
  );
  delay_229 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_349_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_229_q_net
  );
  delay_23 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_156_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_23_q_net
  );
  delay_230 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_350_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_230_q_net
  );
  delay_231 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_351_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_231_q_net
  );
  delay_232 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_352_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_232_q_net
  );
  delay_233 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_353_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_233_q_net
  );
  delay_234 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_354_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_234_q_net
  );
  delay_235 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_355_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_235_q_net
  );
  delay_236 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_356_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_236_q_net
  );
  delay_237 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_357_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_237_q_net
  );
  delay_238 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_358_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_238_q_net
  );
  delay_239 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_359_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_239_q_net
  );
  delay_24 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_157_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_24_q_net
  );
  delay_240 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_360_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_240_q_net
  );
  delay_241 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_361_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_241_q_net
  );
  delay_242 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_362_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_242_q_net
  );
  delay_243 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_363_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_243_q_net
  );
  delay_244 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_364_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_244_q_net
  );
  delay_245 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_365_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_245_q_net
  );
  delay_246 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_366_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_246_q_net
  );
  delay_247 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_367_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_247_q_net
  );
  delay_248 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_368_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_248_q_net
  );
  delay_249 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_369_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_249_q_net
  );
  delay_25 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_158_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_25_q_net
  );
  delay_250 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_370_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_250_q_net
  );
  delay_251 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_371_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_251_q_net
  );
  delay_252 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_372_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_252_q_net
  );
  delay_253 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_373_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_253_q_net
  );
  delay_254 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_374_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_254_q_net
  );
  delay_255 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_375_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_255_q_net
  );
  delay_256 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_376_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_256_q_net
  );
  delay_257 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_377_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_257_q_net
  );
  delay_258 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_378_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_258_q_net
  );
  delay_259 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_379_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_259_q_net
  );
  delay_26 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_159_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_26_q_net
  );
  delay_260 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_380_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_260_q_net
  );
  delay_261 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_381_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_261_q_net
  );
  delay_262 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_382_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_262_q_net
  );
  delay_263 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_383_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_263_q_net
  );
  delay_264 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_384_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_264_q_net
  );
  delay_265 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_385_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_265_q_net
  );
  delay_266 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_386_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_266_q_net
  );
  delay_267 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_387_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_267_q_net
  );
  delay_268 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_388_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_268_q_net
  );
  delay_269 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_389_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_269_q_net
  );
  delay_27 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_160_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_27_q_net
  );
  delay_270 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_390_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_270_q_net
  );
  delay_271 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_391_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_271_q_net
  );
  delay_272 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_392_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_272_q_net
  );
  delay_273 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_393_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_273_q_net
  );
  delay_274 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_394_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_274_q_net
  );
  delay_275 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_395_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_275_q_net
  );
  delay_276 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_396_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_276_q_net
  );
  delay_277 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_397_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_277_q_net
  );
  delay_278 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_398_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_278_q_net
  );
  delay_279 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_399_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_279_q_net
  );
  delay_28 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_161_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_28_q_net
  );
  delay_280 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_400_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_280_q_net
  );
  delay_281 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_401_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_281_q_net
  );
  delay_282 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_402_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_282_q_net
  );
  delay_283 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_403_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_283_q_net
  );
  delay_284 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_404_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_284_q_net
  );
  delay_285 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_405_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_285_q_net
  );
  delay_286 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_406_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_286_q_net
  );
  delay_287 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_407_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_287_q_net
  );
  delay_288 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_408_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_288_q_net
  );
  delay_289 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_409_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_289_q_net
  );
  delay_29 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_162_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_29_q_net
  );
  delay_290 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_410_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_290_q_net
  );
  delay_291 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_411_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_291_q_net
  );
  delay_292 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_412_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_292_q_net
  );
  delay_293 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_413_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_293_q_net
  );
  delay_294 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_414_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_294_q_net
  );
  delay_295 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_415_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_295_q_net
  );
  delay_296 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_416_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_296_q_net
  );
  delay_297 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_417_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_297_q_net
  );
  delay_298 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_418_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_298_q_net
  );
  delay_299 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_419_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_299_q_net
  );
  delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_163_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_3_q_net
  );
  delay_30 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_164_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_30_q_net
  );
  delay_300 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_420_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_300_q_net
  );
  delay_301 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_421_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_301_q_net
  );
  delay_302 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_422_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_302_q_net
  );
  delay_303 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_423_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_303_q_net
  );
  delay_304 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_424_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_304_q_net
  );
  delay_305 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_425_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_305_q_net
  );
  delay_306 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_426_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_306_q_net
  );
  delay_307 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_427_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_307_q_net
  );
  delay_308 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_428_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_308_q_net
  );
  delay_309 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_429_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_309_q_net
  );
  delay_31 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_165_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_31_q_net
  );
  delay_310 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_430_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_310_q_net
  );
  delay_311 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_431_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_311_q_net
  );
  delay_312 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_432_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_312_q_net
  );
  delay_313 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_433_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_313_q_net
  );
  delay_314 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_434_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_314_q_net
  );
  delay_315 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_435_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_315_q_net
  );
  delay_316 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_436_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_316_q_net
  );
  delay_317 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_437_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_317_q_net
  );
  delay_318 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_438_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_318_q_net
  );
  delay_319 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_439_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_319_q_net
  );
  delay_32 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_166_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_32_q_net
  );
  delay_320 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_440_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_320_q_net
  );
  delay_321 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_441_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_321_q_net
  );
  delay_322 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_442_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_322_q_net
  );
  delay_323 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_443_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_323_q_net
  );
  delay_324 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_444_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_324_q_net
  );
  delay_325 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_445_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_325_q_net
  );
  delay_326 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_446_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_326_q_net
  );
  delay_327 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_447_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_327_q_net
  );
  delay_328 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_448_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_328_q_net
  );
  delay_329 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_449_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_329_q_net
  );
  delay_33 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_167_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_33_q_net
  );
  delay_330 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_450_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_330_q_net
  );
  delay_331 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_451_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_331_q_net
  );
  delay_332 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_452_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_332_q_net
  );
  delay_333 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_453_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_333_q_net
  );
  delay_334 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_454_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_334_q_net
  );
  delay_335 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_455_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_335_q_net
  );
  delay_336 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_456_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_336_q_net
  );
  delay_337 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_457_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_337_q_net
  );
  delay_338 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_458_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_338_q_net
  );
  delay_339 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_459_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_339_q_net
  );
  delay_34 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_168_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_34_q_net
  );
  delay_340 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_460_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_340_q_net
  );
  delay_341 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_461_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_341_q_net
  );
  delay_342 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_462_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_342_q_net
  );
  delay_343 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_463_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_343_q_net
  );
  delay_344 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_464_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_344_q_net
  );
  delay_345 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_465_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_345_q_net
  );
  delay_346 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_466_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_346_q_net
  );
  delay_347 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_467_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_347_q_net
  );
  delay_348 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_468_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_348_q_net
  );
  delay_349 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_469_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_349_q_net
  );
  delay_35 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_169_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_35_q_net
  );
  delay_350 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_470_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_350_q_net
  );
  delay_351 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_471_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_351_q_net
  );
  delay_352 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_472_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_352_q_net
  );
  delay_353 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_473_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_353_q_net
  );
  delay_354 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_474_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_354_q_net
  );
  delay_355 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_475_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_355_q_net
  );
  delay_356 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_476_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_356_q_net
  );
  delay_357 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_477_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_357_q_net
  );
  delay_358 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_478_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_358_q_net
  );
  delay_359 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_479_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_359_q_net
  );
  delay_36 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_170_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_36_q_net
  );
  delay_360 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_480_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_360_q_net
  );
  delay_361 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_481_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_361_q_net
  );
  delay_362 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_482_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_362_q_net
  );
  delay_363 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_483_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_363_q_net
  );
  delay_364 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_484_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_364_q_net
  );
  delay_365 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_485_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_365_q_net
  );
  delay_366 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_486_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_366_q_net
  );
  delay_367 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_487_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_367_q_net
  );
  delay_368 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_488_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_368_q_net
  );
  delay_369 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_489_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_369_q_net
  );
  delay_37 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_171_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_37_q_net
  );
  delay_370 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_490_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_370_q_net
  );
  delay_371 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_491_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_371_q_net
  );
  delay_372 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_492_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_372_q_net
  );
  delay_373 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_493_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_373_q_net
  );
  delay_374 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_494_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_374_q_net
  );
  delay_375 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_495_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_375_q_net
  );
  delay_376 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_496_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_376_q_net
  );
  delay_377 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_497_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_377_q_net
  );
  delay_378 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_498_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_378_q_net
  );
  delay_379 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_499_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_379_q_net
  );
  delay_38 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_172_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_38_q_net
  );
  delay_380 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_500_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_380_q_net
  );
  delay_381 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_501_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_381_q_net
  );
  delay_382 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_502_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_382_q_net
  );
  delay_383 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_503_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_383_q_net
  );
  delay_384 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_504_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_384_q_net
  );
  delay_385 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_505_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_385_q_net
  );
  delay_386 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_506_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_386_q_net
  );
  delay_387 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_507_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_387_q_net
  );
  delay_388 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_508_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_388_q_net
  );
  delay_389 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_509_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_389_q_net
  );
  delay_39 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_173_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_39_q_net
  );
  delay_390 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_510_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_390_q_net
  );
  delay_391 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_511_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_391_q_net
  );
  delay_392 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_512_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_392_q_net
  );
  delay_393 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_513_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_393_q_net
  );
  delay_394 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_514_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_394_q_net
  );
  delay_395 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_515_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_395_q_net
  );
  delay_396 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_516_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_396_q_net
  );
  delay_397 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_517_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_397_q_net
  );
  delay_398 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_518_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_398_q_net
  );
  delay_399 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_519_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_399_q_net
  );
  delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_174_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_4_q_net
  );
  delay_40 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_175_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_40_q_net
  );
  delay_400 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_520_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_400_q_net
  );
  delay_401 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_521_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_401_q_net
  );
  delay_402 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_522_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_402_q_net
  );
  delay_403 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_523_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_403_q_net
  );
  delay_404 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_524_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_404_q_net
  );
  delay_405 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_525_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_405_q_net
  );
  delay_406 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_526_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_406_q_net
  );
  delay_407 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_527_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_407_q_net
  );
  delay_408 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_528_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_408_q_net
  );
  delay_409 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_529_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_409_q_net
  );
  delay_41 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_176_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_41_q_net
  );
  delay_410 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_530_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_410_q_net
  );
  delay_411 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_531_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_411_q_net
  );
  delay_412 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_532_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_412_q_net
  );
  delay_413 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_533_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_413_q_net
  );
  delay_414 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_534_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_414_q_net
  );
  delay_415 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_535_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_415_q_net
  );
  delay_416 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_536_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_416_q_net
  );
  delay_417 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_537_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_417_q_net
  );
  delay_418 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_538_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_418_q_net
  );
  delay_419 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_539_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_419_q_net
  );
  delay_42 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_177_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_42_q_net
  );
  delay_420 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_540_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_420_q_net
  );
  delay_421 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_541_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_421_q_net
  );
  delay_422 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_542_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_422_q_net
  );
  delay_423 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_543_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_423_q_net
  );
  delay_424 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_544_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_424_q_net
  );
  delay_425 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_545_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_425_q_net
  );
  delay_426 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_546_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_426_q_net
  );
  delay_427 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_547_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_427_q_net
  );
  delay_428 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_548_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_428_q_net
  );
  delay_429 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_549_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_429_q_net
  );
  delay_43 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_178_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_43_q_net
  );
  delay_430 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_550_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_430_q_net
  );
  delay_431 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_551_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_431_q_net
  );
  delay_432 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_552_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_432_q_net
  );
  delay_433 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_553_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_433_q_net
  );
  delay_434 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_554_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_434_q_net
  );
  delay_435 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_555_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_435_q_net
  );
  delay_436 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_556_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_436_q_net
  );
  delay_437 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_557_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_437_q_net
  );
  delay_438 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_558_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_438_q_net
  );
  delay_439 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_559_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_439_q_net
  );
  delay_44 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_179_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_44_q_net
  );
  delay_440 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_560_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_440_q_net
  );
  delay_441 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_561_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_441_q_net
  );
  delay_442 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_562_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_442_q_net
  );
  delay_443 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_563_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_443_q_net
  );
  delay_444 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_564_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_444_q_net
  );
  delay_445 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_565_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_445_q_net
  );
  delay_446 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_566_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_446_q_net
  );
  delay_447 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_567_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_447_q_net
  );
  delay_448 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_568_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_448_q_net
  );
  delay_449 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_569_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_449_q_net
  );
  delay_45 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_180_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_45_q_net
  );
  delay_450 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_570_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_450_q_net
  );
  delay_451 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_571_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_451_q_net
  );
  delay_452 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_572_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_452_q_net
  );
  delay_453 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_573_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_453_q_net
  );
  delay_454 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_574_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_454_q_net
  );
  delay_455 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_575_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_455_q_net
  );
  delay_456 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_576_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_456_q_net
  );
  delay_457 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_577_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_457_q_net
  );
  delay_458 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_578_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_458_q_net
  );
  delay_459 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_579_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_459_q_net
  );
  delay_46 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_181_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_46_q_net
  );
  delay_460 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_580_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_460_q_net
  );
  delay_461 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_581_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_461_q_net
  );
  delay_462 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_582_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_462_q_net
  );
  delay_463 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_583_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_463_q_net
  );
  delay_464 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_584_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_464_q_net
  );
  delay_465 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_585_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_465_q_net
  );
  delay_466 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_586_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_466_q_net
  );
  delay_467 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_587_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_467_q_net
  );
  delay_468 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_588_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_468_q_net
  );
  delay_469 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_589_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_469_q_net
  );
  delay_47 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_182_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_47_q_net
  );
  delay_470 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_590_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_470_q_net
  );
  delay_471 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_591_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_471_q_net
  );
  delay_472 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_592_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_472_q_net
  );
  delay_473 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_593_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_473_q_net
  );
  delay_474 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_594_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_474_q_net
  );
  delay_475 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_595_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_475_q_net
  );
  delay_476 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_596_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_476_q_net
  );
  delay_477 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_597_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_477_q_net
  );
  delay_478 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_598_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_478_q_net
  );
  delay_479 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_599_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_479_q_net
  );
  delay_48 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_183_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_48_q_net
  );
  delay_480 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_600_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_480_q_net
  );
  delay_481 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_601_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_481_q_net
  );
  delay_482 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_602_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_482_q_net
  );
  delay_483 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_603_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_483_q_net
  );
  delay_484 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_604_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_484_q_net
  );
  delay_485 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_605_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_485_q_net
  );
  delay_486 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_606_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_486_q_net
  );
  delay_487 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_607_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_487_q_net
  );
  delay_488 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_608_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_488_q_net
  );
  delay_489 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_609_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_489_q_net
  );
  delay_49 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_184_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_49_q_net
  );
  delay_490 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_610_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_490_q_net
  );
  delay_491 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_611_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_491_q_net
  );
  delay_492 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_612_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_492_q_net
  );
  delay_493 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_613_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_493_q_net
  );
  delay_494 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_614_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_494_q_net
  );
  delay_495 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_615_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_495_q_net
  );
  delay_496 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_616_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_496_q_net
  );
  delay_497 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_617_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_497_q_net
  );
  delay_498 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_618_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_498_q_net
  );
  delay_499 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_619_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_499_q_net
  );
  delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_185_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_5_q_net
  );
  delay_50 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_186_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_50_q_net
  );
  delay_500 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_620_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_500_q_net
  );
  delay_501 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_621_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_501_q_net
  );
  delay_502 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_622_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_502_q_net
  );
  delay_503 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_623_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_503_q_net
  );
  delay_504 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_624_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_504_q_net
  );
  delay_505 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_625_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_505_q_net
  );
  delay_506 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_626_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_506_q_net
  );
  delay_507 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_627_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_507_q_net
  );
  delay_508 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_628_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_508_q_net
  );
  delay_509 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_629_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_509_q_net
  );
  delay_51 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_187_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_51_q_net
  );
  delay_510 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_630_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_510_q_net
  );
  delay_511 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_631_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_511_q_net
  );
  delay_512 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_632_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_512_q_net
  );
  delay_513 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_633_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_513_q_net
  );
  delay_514 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_634_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_514_q_net
  );
  delay_515 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_635_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_515_q_net
  );
  delay_516 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_636_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_516_q_net
  );
  delay_517 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_637_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_517_q_net
  );
  delay_518 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_638_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_518_q_net
  );
  delay_519 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_639_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_519_q_net
  );
  delay_52 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_188_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_52_q_net
  );
  delay_520 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_640_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_520_q_net
  );
  delay_521 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_641_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_521_q_net
  );
  delay_522 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_642_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_522_q_net
  );
  delay_523 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_643_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_523_q_net
  );
  delay_524 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_644_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_524_q_net
  );
  delay_525 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_645_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_525_q_net
  );
  delay_526 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_646_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_526_q_net
  );
  delay_527 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_647_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_527_q_net
  );
  delay_528 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_648_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_528_q_net
  );
  delay_529 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_649_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_529_q_net
  );
  delay_53 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_189_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_53_q_net
  );
  delay_530 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_650_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_530_q_net
  );
  delay_531 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_651_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_531_q_net
  );
  delay_532 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_652_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_532_q_net
  );
  delay_533 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_653_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_533_q_net
  );
  delay_534 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_654_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_534_q_net
  );
  delay_535 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_655_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_535_q_net
  );
  delay_536 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_656_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_536_q_net
  );
  delay_537 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_657_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_537_q_net
  );
  delay_538 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_658_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_538_q_net
  );
  delay_539 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_659_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_539_q_net
  );
  delay_54 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_190_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_54_q_net
  );
  delay_540 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_660_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_540_q_net
  );
  delay_541 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_661_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_541_q_net
  );
  delay_542 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_662_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_542_q_net
  );
  delay_543 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_663_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_543_q_net
  );
  delay_544 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_664_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_544_q_net
  );
  delay_545 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_665_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_545_q_net
  );
  delay_546 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_666_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_546_q_net
  );
  delay_547 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_667_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_547_q_net
  );
  delay_548 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_668_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_548_q_net
  );
  delay_549 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_669_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_549_q_net
  );
  delay_55 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_191_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_55_q_net
  );
  delay_550 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_670_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_550_q_net
  );
  delay_551 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_671_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_551_q_net
  );
  delay_552 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_672_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_552_q_net
  );
  delay_553 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_673_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_553_q_net
  );
  delay_554 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_674_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_554_q_net
  );
  delay_555 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_675_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_555_q_net
  );
  delay_556 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_676_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_556_q_net
  );
  delay_557 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_677_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_557_q_net
  );
  delay_558 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_678_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_558_q_net
  );
  delay_559 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_679_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_559_q_net
  );
  delay_56 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_192_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_56_q_net
  );
  delay_560 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_680_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_560_q_net
  );
  delay_561 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_681_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_561_q_net
  );
  delay_562 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_682_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_562_q_net
  );
  delay_563 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_683_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_563_q_net
  );
  delay_564 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_684_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_564_q_net
  );
  delay_565 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_685_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_565_q_net
  );
  delay_566 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_686_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_566_q_net
  );
  delay_567 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_687_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_567_q_net
  );
  delay_568 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_688_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_568_q_net
  );
  delay_569 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_689_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_569_q_net
  );
  delay_57 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_193_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_57_q_net
  );
  delay_570 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_690_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_570_q_net
  );
  delay_571 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_691_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_571_q_net
  );
  delay_572 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_692_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_572_q_net
  );
  delay_573 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_693_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_573_q_net
  );
  delay_574 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_694_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_574_q_net
  );
  delay_575 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_695_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_575_q_net
  );
  delay_576 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_696_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_576_q_net
  );
  delay_577 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_697_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_577_q_net
  );
  delay_578 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_698_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_578_q_net
  );
  delay_579 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_699_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_579_q_net
  );
  delay_58 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_194_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_58_q_net
  );
  delay_580 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_700_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_580_q_net
  );
  delay_581 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_701_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_581_q_net
  );
  delay_582 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_702_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_582_q_net
  );
  delay_583 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_703_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_583_q_net
  );
  delay_584 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_704_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_584_q_net
  );
  delay_585 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_705_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_585_q_net
  );
  delay_586 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_706_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_586_q_net
  );
  delay_587 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_707_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_587_q_net
  );
  delay_588 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_708_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_588_q_net
  );
  delay_589 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_709_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_589_q_net
  );
  delay_59 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_195_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_59_q_net
  );
  delay_590 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_710_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_590_q_net
  );
  delay_591 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_711_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_591_q_net
  );
  delay_592 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_712_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_592_q_net
  );
  delay_593 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_713_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_593_q_net
  );
  delay_594 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_714_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_594_q_net
  );
  delay_595 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_715_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_595_q_net
  );
  delay_596 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_716_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_596_q_net
  );
  delay_597 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_717_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_597_q_net
  );
  delay_598 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_718_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_598_q_net
  );
  delay_599 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_719_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_599_q_net
  );
  delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_196_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_6_q_net
  );
  delay_60 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_197_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_60_q_net
  );
  delay_600 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_840_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_600_q_net
  );
  delay_601 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_841_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_601_q_net
  );
  delay_602 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_842_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_602_q_net
  );
  delay_603 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_843_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_603_q_net
  );
  delay_604 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_844_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_604_q_net
  );
  delay_605 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_845_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_605_q_net
  );
  delay_606 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_846_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_606_q_net
  );
  delay_607 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_847_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_607_q_net
  );
  delay_608 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_848_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_608_q_net
  );
  delay_609 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_849_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_609_q_net
  );
  delay_61 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_198_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_61_q_net
  );
  delay_610 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_850_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_610_q_net
  );
  delay_611 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_851_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_611_q_net
  );
  delay_612 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_852_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_612_q_net
  );
  delay_613 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_853_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_613_q_net
  );
  delay_614 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_854_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_614_q_net
  );
  delay_615 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_855_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_615_q_net
  );
  delay_616 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_856_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_616_q_net
  );
  delay_617 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_857_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_617_q_net
  );
  delay_618 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_858_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_618_q_net
  );
  delay_619 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_859_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_619_q_net
  );
  delay_62 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_199_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_62_q_net
  );
  delay_620 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_860_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_620_q_net
  );
  delay_621 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_861_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_621_q_net
  );
  delay_622 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_862_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_622_q_net
  );
  delay_623 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_863_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_623_q_net
  );
  delay_624 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_864_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_624_q_net
  );
  delay_625 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_865_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_625_q_net
  );
  delay_626 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_866_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_626_q_net
  );
  delay_627 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_867_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_627_q_net
  );
  delay_628 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_868_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_628_q_net
  );
  delay_629 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_869_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_629_q_net
  );
  delay_63 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_200_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_63_q_net
  );
  delay_630 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_870_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_630_q_net
  );
  delay_631 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_871_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_631_q_net
  );
  delay_632 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_872_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_632_q_net
  );
  delay_633 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_873_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_633_q_net
  );
  delay_634 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_874_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_634_q_net
  );
  delay_635 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_875_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_635_q_net
  );
  delay_636 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_876_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_636_q_net
  );
  delay_637 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_877_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_637_q_net
  );
  delay_638 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_878_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_638_q_net
  );
  delay_639 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_879_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_639_q_net
  );
  delay_64 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_201_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_64_q_net
  );
  delay_640 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_880_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_640_q_net
  );
  delay_641 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_881_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_641_q_net
  );
  delay_642 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_882_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_642_q_net
  );
  delay_643 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_883_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_643_q_net
  );
  delay_644 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_884_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_644_q_net
  );
  delay_645 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_885_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_645_q_net
  );
  delay_646 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_886_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_646_q_net
  );
  delay_647 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_887_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_647_q_net
  );
  delay_648 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_888_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_648_q_net
  );
  delay_649 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_889_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_649_q_net
  );
  delay_65 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_202_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_65_q_net
  );
  delay_650 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_890_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_650_q_net
  );
  delay_651 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_891_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_651_q_net
  );
  delay_652 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_892_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_652_q_net
  );
  delay_653 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_893_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_653_q_net
  );
  delay_654 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_894_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_654_q_net
  );
  delay_655 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_895_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_655_q_net
  );
  delay_656 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_896_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_656_q_net
  );
  delay_657 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_897_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_657_q_net
  );
  delay_658 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_898_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_658_q_net
  );
  delay_659 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_899_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_659_q_net
  );
  delay_66 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_203_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_66_q_net
  );
  delay_660 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_900_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_660_q_net
  );
  delay_661 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_901_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_661_q_net
  );
  delay_662 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_902_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_662_q_net
  );
  delay_663 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_903_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_663_q_net
  );
  delay_664 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_904_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_664_q_net
  );
  delay_665 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_905_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_665_q_net
  );
  delay_666 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_906_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_666_q_net
  );
  delay_667 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_907_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_667_q_net
  );
  delay_668 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_908_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_668_q_net
  );
  delay_669 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_909_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_669_q_net
  );
  delay_67 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_204_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_67_q_net
  );
  delay_670 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_910_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_670_q_net
  );
  delay_671 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_911_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_671_q_net
  );
  delay_672 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_912_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_672_q_net
  );
  delay_673 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_913_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_673_q_net
  );
  delay_674 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_914_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_674_q_net
  );
  delay_675 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_915_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_675_q_net
  );
  delay_676 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_916_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_676_q_net
  );
  delay_677 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_917_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_677_q_net
  );
  delay_678 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_918_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_678_q_net
  );
  delay_679 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_919_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_679_q_net
  );
  delay_68 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_205_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_68_q_net
  );
  delay_680 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_920_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_680_q_net
  );
  delay_681 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_921_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_681_q_net
  );
  delay_682 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_922_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_682_q_net
  );
  delay_683 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_923_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_683_q_net
  );
  delay_684 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_924_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_684_q_net
  );
  delay_685 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_925_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_685_q_net
  );
  delay_686 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_926_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_686_q_net
  );
  delay_687 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_927_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_687_q_net
  );
  delay_688 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_928_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_688_q_net
  );
  delay_689 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_929_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_689_q_net
  );
  delay_69 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_206_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_69_q_net
  );
  delay_690 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_930_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_690_q_net
  );
  delay_691 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_931_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_691_q_net
  );
  delay_692 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_932_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_692_q_net
  );
  delay_693 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_933_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_693_q_net
  );
  delay_694 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_934_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_694_q_net
  );
  delay_695 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_935_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_695_q_net
  );
  delay_696 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_936_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_696_q_net
  );
  delay_697 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_937_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_697_q_net
  );
  delay_698 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_938_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_698_q_net
  );
  delay_699 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_939_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_699_q_net
  );
  delay_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_207_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_7_q_net
  );
  delay_70 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_208_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_70_q_net
  );
  delay_700 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_940_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_700_q_net
  );
  delay_701 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_941_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_701_q_net
  );
  delay_702 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_942_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_702_q_net
  );
  delay_703 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_943_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_703_q_net
  );
  delay_704 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_944_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_704_q_net
  );
  delay_705 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_945_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_705_q_net
  );
  delay_706 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_946_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_706_q_net
  );
  delay_707 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_947_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_707_q_net
  );
  delay_708 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_948_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_708_q_net
  );
  delay_709 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_949_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_709_q_net
  );
  delay_71 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_209_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_71_q_net
  );
  delay_710 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_950_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_710_q_net
  );
  delay_711 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_951_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_711_q_net
  );
  delay_712 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_952_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_712_q_net
  );
  delay_713 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_953_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_713_q_net
  );
  delay_714 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_954_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_714_q_net
  );
  delay_715 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_955_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_715_q_net
  );
  delay_716 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_956_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_716_q_net
  );
  delay_717 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_957_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_717_q_net
  );
  delay_718 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_958_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_718_q_net
  );
  delay_719 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_959_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_719_q_net
  );
  delay_72 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_210_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_72_q_net
  );
  delay_720 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_720_q_net
  );
  delay_721 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_721_q_net
  );
  delay_722 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_722_q_net
  );
  delay_723 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_723_q_net
  );
  delay_724 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_724_q_net
  );
  delay_725 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_725_q_net
  );
  delay_726 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_726_q_net
  );
  delay_727 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_727_q_net
  );
  delay_728 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_728_q_net
  );
  delay_729 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_729_q_net
  );
  delay_73 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_211_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_73_q_net
  );
  delay_730 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_730_q_net
  );
  delay_731 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_731_q_net
  );
  delay_732 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_732_q_net
  );
  delay_733 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_733_q_net
  );
  delay_734 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_734_q_net
  );
  delay_735 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_735_q_net
  );
  delay_736 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_736_q_net
  );
  delay_737 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_737_q_net
  );
  delay_738 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_738_q_net
  );
  delay_739 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_739_q_net
  );
  delay_74 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_212_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_74_q_net
  );
  delay_740 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_740_q_net
  );
  delay_741 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_741_q_net
  );
  delay_742 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_742_q_net
  );
  delay_743 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_743_q_net
  );
  delay_744 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_744_q_net
  );
  delay_745 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_745_q_net
  );
  delay_746 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_746_q_net
  );
  delay_747 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_747_q_net
  );
  delay_748 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_748_q_net
  );
  delay_749 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_749_q_net
  );
  delay_75 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_213_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_75_q_net
  );
  delay_750 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_750_q_net
  );
  delay_751 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_751_q_net
  );
  delay_752 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_752_q_net
  );
  delay_753 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_753_q_net
  );
  delay_754 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_754_q_net
  );
  delay_755 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_755_q_net
  );
  delay_756 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_756_q_net
  );
  delay_757 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_757_q_net
  );
  delay_758 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_758_q_net
  );
  delay_759 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_759_q_net
  );
  delay_76 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_214_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_76_q_net
  );
  delay_760 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_760_q_net
  );
  delay_761 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_761_q_net
  );
  delay_762 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_762_q_net
  );
  delay_763 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_763_q_net
  );
  delay_764 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_764_q_net
  );
  delay_765 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_765_q_net
  );
  delay_766 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_766_q_net
  );
  delay_767 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_767_q_net
  );
  delay_768 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_768_q_net
  );
  delay_769 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_769_q_net
  );
  delay_77 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_215_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_77_q_net
  );
  delay_770 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_770_q_net
  );
  delay_771 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_771_q_net
  );
  delay_772 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_772_q_net
  );
  delay_773 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_773_q_net
  );
  delay_774 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_774_q_net
  );
  delay_775 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_775_q_net
  );
  delay_776 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_776_q_net
  );
  delay_777 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_777_q_net
  );
  delay_778 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_778_q_net
  );
  delay_779 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_779_q_net
  );
  delay_78 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_216_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_78_q_net
  );
  delay_780 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_780_q_net
  );
  delay_781 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay_781_q_net
  );
  delay_782 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_782_q_net
  );
  delay_783 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_783_q_net
  );
  delay_784 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_784_q_net
  );
  delay_785 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_785_q_net
  );
  delay_786 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_786_q_net
  );
  delay_787 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_787_q_net
  );
  delay_788 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_788_q_net
  );
  delay_789 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_789_q_net
  );
  delay_79 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_217_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_79_q_net
  );
  delay_790 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_790_q_net
  );
  delay_791 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_791_q_net
  );
  delay_792 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_792_q_net
  );
  delay_793 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_793_q_net
  );
  delay_794 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_794_q_net
  );
  delay_795 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_795_q_net
  );
  delay_796 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_796_q_net
  );
  delay_797 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_797_q_net
  );
  delay_798 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_798_q_net
  );
  delay_799 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_799_q_net
  );
  delay_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_218_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_8_q_net
  );
  delay_80 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_219_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_80_q_net
  );
  delay_800 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_800_q_net
  );
  delay_801 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_801_q_net
  );
  delay_802 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_802_q_net
  );
  delay_803 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_803_q_net
  );
  delay_804 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_804_q_net
  );
  delay_805 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_805_q_net
  );
  delay_806 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_806_q_net
  );
  delay_807 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_807_q_net
  );
  delay_808 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay_808_q_net
  );
  delay_809 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay_809_q_net
  );
  delay_81 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_220_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_81_q_net
  );
  delay_810 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_810_q_net
  );
  delay_811 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_811_q_net
  );
  delay_812 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_812_q_net
  );
  delay_813 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_813_q_net
  );
  delay_814 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_814_q_net
  );
  delay_815 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_815_q_net
  );
  delay_816 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_816_q_net
  );
  delay_817 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_7_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_817_q_net
  );
  delay_818 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_818_q_net
  );
  delay_819 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_819_q_net
  );
  delay_82 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_221_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_82_q_net
  );
  delay_820 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_9_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_820_q_net
  );
  delay_821 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_821_q_net
  );
  delay_822 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_10_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_822_q_net
  );
  delay_823 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_823_q_net
  );
  delay_824 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_824_q_net
  );
  delay_825 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_11_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_825_q_net
  );
  delay_826 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_826_q_net
  );
  delay_827 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_8_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_827_q_net
  );
  delay_828 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_1_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_828_q_net
  );
  delay_829 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay_829_q_net
  );
  delay_83 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_222_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_83_q_net
  );
  delay_830 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_830_q_net
  );
  delay_831 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_2_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_831_q_net
  );
  delay_832 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_832_q_net
  );
  delay_833 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_3_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_833_q_net
  );
  delay_834 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay_834_q_net
  );
  delay_835 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_835_q_net
  );
  delay_836 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_836_q_net
  );
  delay_837 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_837_q_net
  );
  delay_838 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay_838_q_net
  );
  delay_839 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => x12_bit_bin_value_5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_839_q_net
  );
  delay_84 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_223_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_84_q_net
  );
  delay_840 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_720_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_840_q_net
  );
  delay_841 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_721_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_841_q_net
  );
  delay_842 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_722_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_842_q_net
  );
  delay_843 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_723_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_843_q_net
  );
  delay_844 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_724_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_844_q_net
  );
  delay_845 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_725_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_845_q_net
  );
  delay_846 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_726_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_846_q_net
  );
  delay_847 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_727_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_847_q_net
  );
  delay_848 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_728_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_848_q_net
  );
  delay_849 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_729_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_849_q_net
  );
  delay_85 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_224_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_85_q_net
  );
  delay_850 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_730_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_850_q_net
  );
  delay_851 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_731_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_851_q_net
  );
  delay_852 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_732_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_852_q_net
  );
  delay_853 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_733_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_853_q_net
  );
  delay_854 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_734_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_854_q_net
  );
  delay_855 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_735_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_855_q_net
  );
  delay_856 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_736_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_856_q_net
  );
  delay_857 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_737_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_857_q_net
  );
  delay_858 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_738_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_858_q_net
  );
  delay_859 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_739_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_859_q_net
  );
  delay_86 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_225_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_86_q_net
  );
  delay_860 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_740_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_860_q_net
  );
  delay_861 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_741_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_861_q_net
  );
  delay_862 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_742_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_862_q_net
  );
  delay_863 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_743_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_863_q_net
  );
  delay_864 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_744_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_864_q_net
  );
  delay_865 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_745_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_865_q_net
  );
  delay_866 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_746_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_866_q_net
  );
  delay_867 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_747_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_867_q_net
  );
  delay_868 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_748_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_868_q_net
  );
  delay_869 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_749_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_869_q_net
  );
  delay_87 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_226_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_87_q_net
  );
  delay_870 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_750_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_870_q_net
  );
  delay_871 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_751_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_871_q_net
  );
  delay_872 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_752_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_872_q_net
  );
  delay_873 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_753_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_873_q_net
  );
  delay_874 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_754_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_874_q_net
  );
  delay_875 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_755_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_875_q_net
  );
  delay_876 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_756_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_876_q_net
  );
  delay_877 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_757_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_877_q_net
  );
  delay_878 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_758_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_878_q_net
  );
  delay_879 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_759_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_879_q_net
  );
  delay_88 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_227_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_88_q_net
  );
  delay_880 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_760_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_880_q_net
  );
  delay_881 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_761_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_881_q_net
  );
  delay_882 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_762_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_882_q_net
  );
  delay_883 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_763_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_883_q_net
  );
  delay_884 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_764_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_884_q_net
  );
  delay_885 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_765_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_885_q_net
  );
  delay_886 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_766_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_886_q_net
  );
  delay_887 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_767_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_887_q_net
  );
  delay_888 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_768_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_888_q_net
  );
  delay_889 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_769_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_889_q_net
  );
  delay_89 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_228_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_89_q_net
  );
  delay_890 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_770_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_890_q_net
  );
  delay_891 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_771_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_891_q_net
  );
  delay_892 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_772_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_892_q_net
  );
  delay_893 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_773_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_893_q_net
  );
  delay_894 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_774_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_894_q_net
  );
  delay_895 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_775_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_895_q_net
  );
  delay_896 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_776_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_896_q_net
  );
  delay_897 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_777_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_897_q_net
  );
  delay_898 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_778_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_898_q_net
  );
  delay_899 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_779_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_899_q_net
  );
  delay_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_229_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_9_q_net
  );
  delay_90 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_230_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_90_q_net
  );
  delay_900 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_780_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_900_q_net
  );
  delay_901 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_781_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_901_q_net
  );
  delay_902 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_782_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_902_q_net
  );
  delay_903 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_783_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_903_q_net
  );
  delay_904 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_784_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_904_q_net
  );
  delay_905 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_785_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_905_q_net
  );
  delay_906 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_786_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_906_q_net
  );
  delay_907 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_787_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_907_q_net
  );
  delay_908 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_788_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_908_q_net
  );
  delay_909 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_789_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_909_q_net
  );
  delay_91 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_231_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_91_q_net
  );
  delay_910 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_790_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_910_q_net
  );
  delay_911 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_791_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_911_q_net
  );
  delay_912 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_792_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_912_q_net
  );
  delay_913 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_793_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_913_q_net
  );
  delay_914 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_794_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_914_q_net
  );
  delay_915 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_795_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_915_q_net
  );
  delay_916 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_796_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_916_q_net
  );
  delay_917 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_797_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_917_q_net
  );
  delay_918 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_798_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_918_q_net
  );
  delay_919 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_799_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_919_q_net
  );
  delay_92 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_232_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_92_q_net
  );
  delay_920 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_800_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_920_q_net
  );
  delay_921 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_801_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_921_q_net
  );
  delay_922 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_802_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_922_q_net
  );
  delay_923 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_803_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_923_q_net
  );
  delay_924 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_804_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_924_q_net
  );
  delay_925 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_805_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_925_q_net
  );
  delay_926 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_806_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_926_q_net
  );
  delay_927 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_807_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_927_q_net
  );
  delay_928 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_808_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_928_q_net
  );
  delay_929 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_809_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_929_q_net
  );
  delay_93 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_233_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_93_q_net
  );
  delay_930 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_810_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_930_q_net
  );
  delay_931 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_811_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_931_q_net
  );
  delay_932 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_812_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_932_q_net
  );
  delay_933 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_813_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_933_q_net
  );
  delay_934 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_814_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_934_q_net
  );
  delay_935 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_815_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_935_q_net
  );
  delay_936 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_816_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_936_q_net
  );
  delay_937 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_817_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_937_q_net
  );
  delay_938 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_818_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_938_q_net
  );
  delay_939 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_819_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_939_q_net
  );
  delay_94 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_234_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_94_q_net
  );
  delay_940 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_820_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_940_q_net
  );
  delay_941 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_821_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_941_q_net
  );
  delay_942 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_822_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_942_q_net
  );
  delay_943 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_823_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_943_q_net
  );
  delay_944 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_824_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_944_q_net
  );
  delay_945 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_825_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_945_q_net
  );
  delay_946 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_826_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_946_q_net
  );
  delay_947 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_827_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_947_q_net
  );
  delay_948 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_828_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_948_q_net
  );
  delay_949 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_829_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_949_q_net
  );
  delay_95 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_235_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_95_q_net
  );
  delay_950 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_830_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_950_q_net
  );
  delay_951 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_831_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_951_q_net
  );
  delay_952 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_832_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_952_q_net
  );
  delay_953 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_833_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_953_q_net
  );
  delay_954 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_834_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_954_q_net
  );
  delay_955 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_835_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_955_q_net
  );
  delay_956 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_836_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_956_q_net
  );
  delay_957 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_837_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_957_q_net
  );
  delay_958 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_838_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_958_q_net
  );
  delay_959 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_839_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_959_q_net
  );
  delay_96 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_236_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_96_q_net
  );
  delay_97 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_237_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_97_q_net
  );
  delay_98 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_238_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_98_q_net
  );
  delay_99 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_239_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_99_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results;
architecture structural of mh_accumlator_kernel_results is 
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0;
architecture structural of mh_accumulator_offset_0 is 
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1;
architecture structural of mh_accumulator_offset_1 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2;
architecture structural of mh_accumulator_offset_2 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3;
architecture structural of mh_accumulator_offset_3 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4;
architecture structural of mh_accumulator_offset_4 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0;
architecture structural of mh_multiple_and_add_offset_0 is 
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1;
architecture structural of mh_multiple_and_add_offset_1 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2;
architecture structural of mh_multiple_and_add_offset_2 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3;
architecture structural of mh_multiple_and_add_offset_3 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4;
architecture structural of mh_multiple_and_add_offset_4 is 
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_0 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_0;
architecture structural of mh_kernel_result_0 is 
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_0_q_net <= pixel_bus_input_offset_0_1;
  delay_22_q_net <= pixel_bus_input_offset_1_1;
  delay_48_q_net <= pixel_bus_input_offset_2_1;
  delay_72_q_net <= pixel_bus_input_offset_3_1;
  delay_96_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_0_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_2_q_net <= pixel_bus_input_offset_0_2;
  delay_4_q_net <= pixel_bus_input_offset_0_3;
  delay_6_q_net <= pixel_bus_input_offset_0_4;
  delay_8_q_net <= pixel_bus_input_offset_0_5;
  delay_10_q_net <= pixel_bus_input_offset_0_6;
  delay_12_q_net <= pixel_bus_input_offset_0_7;
  delay_14_q_net <= pixel_bus_input_offset_0_8;
  delay_23_q_net <= pixel_bus_input_offset_0_9;
  delay_16_q_net <= pixel_bus_input_offset_0_10;
  delay_18_q_net <= pixel_bus_input_offset_0_11;
  delay_20_q_net <= pixel_bus_input_offset_0_12;
  delay_36_q_net <= pixel_bus_input_offset_1_2;
  delay_42_q_net <= pixel_bus_input_offset_1_3;
  delay_44_q_net <= pixel_bus_input_offset_1_4;
  delay_46_q_net <= pixel_bus_input_offset_1_5;
  delay_26_q_net <= pixel_bus_input_offset_1_6;
  delay_28_q_net <= pixel_bus_input_offset_1_7;
  delay_30_q_net <= pixel_bus_input_offset_1_8;
  delay_39_q_net <= pixel_bus_input_offset_1_9;
  delay_32_q_net <= pixel_bus_input_offset_1_10;
  delay_34_q_net <= pixel_bus_input_offset_1_11;
  delay_37_q_net <= pixel_bus_input_offset_1_12;
  delay_60_q_net <= pixel_bus_input_offset_2_2;
  delay_66_q_net <= pixel_bus_input_offset_2_3;
  delay_68_q_net <= pixel_bus_input_offset_2_4;
  delay_70_q_net <= pixel_bus_input_offset_2_5;
  delay_50_q_net <= pixel_bus_input_offset_2_6;
  delay_52_q_net <= pixel_bus_input_offset_2_7;
  delay_54_q_net <= pixel_bus_input_offset_2_8;
  delay_63_q_net <= pixel_bus_input_offset_2_9;
  delay_56_q_net <= pixel_bus_input_offset_2_10;
  delay_58_q_net <= pixel_bus_input_offset_2_11;
  delay_61_q_net <= pixel_bus_input_offset_2_12;
  delay_84_q_net <= pixel_bus_input_offset_3_2;
  delay_90_q_net <= pixel_bus_input_offset_3_3;
  delay_92_q_net <= pixel_bus_input_offset_3_4;
  delay_94_q_net <= pixel_bus_input_offset_3_5;
  delay_74_q_net <= pixel_bus_input_offset_3_6;
  delay_76_q_net <= pixel_bus_input_offset_3_7;
  delay_78_q_net <= pixel_bus_input_offset_3_8;
  delay_87_q_net <= pixel_bus_input_offset_3_9;
  delay_80_q_net <= pixel_bus_input_offset_3_10;
  delay_82_q_net <= pixel_bus_input_offset_3_11;
  delay_85_q_net <= pixel_bus_input_offset_3_12;
  delay_108_q_net <= pixel_bus_input_offset_4_2;
  delay_114_q_net <= pixel_bus_input_offset_4_3;
  delay_116_q_net <= pixel_bus_input_offset_4_4;
  delay_118_q_net <= pixel_bus_input_offset_4_5;
  delay_98_q_net <= pixel_bus_input_offset_4_6;
  delay_100_q_net <= pixel_bus_input_offset_4_7;
  delay_102_q_net <= pixel_bus_input_offset_4_8;
  delay_111_q_net <= pixel_bus_input_offset_4_9;
  delay_104_q_net <= pixel_bus_input_offset_4_10;
  delay_106_q_net <= pixel_bus_input_offset_4_11;
  delay_109_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x0 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x0;
architecture structural of mh_accumlator_kernel_results_x0 is 
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x0 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x0;
architecture structural of mh_accumulator_offset_0_x0 is 
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x0 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x0;
architecture structural of mh_accumulator_offset_1_x0 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x0 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x0;
architecture structural of mh_accumulator_offset_2_x0 is 
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x0 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x0;
architecture structural of mh_accumulator_offset_3_x0 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x0 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x0;
architecture structural of mh_accumulator_offset_4_x0 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x0 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x0;
architecture structural of mh_multiple_and_add_offset_0_x0 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x0 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x0;
architecture structural of mh_multiple_and_add_offset_1_x0 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x0 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x0;
architecture structural of mh_multiple_and_add_offset_2_x0 is 
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x0 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x0;
architecture structural of mh_multiple_and_add_offset_3_x0 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x0 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x0;
architecture structural of mh_multiple_and_add_offset_4_x0 is 
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_1 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_5 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_1;
architecture structural of mh_kernel_result_1 is 
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_22_q_net <= pixel_bus_input_offset_0_1;
  delay_48_q_net <= pixel_bus_input_offset_1_1;
  delay_72_q_net <= pixel_bus_input_offset_2_1;
  delay_96_q_net <= pixel_bus_input_offset_3_1;
  delay_0_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_0_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_36_q_net <= pixel_bus_input_offset_0_2;
  delay_42_q_net <= pixel_bus_input_offset_0_3;
  delay_44_q_net <= pixel_bus_input_offset_0_4;
  delay_46_q_net <= pixel_bus_input_offset_0_5;
  delay_26_q_net <= pixel_bus_input_offset_0_6;
  delay_28_q_net <= pixel_bus_input_offset_0_7;
  delay_30_q_net <= pixel_bus_input_offset_0_8;
  delay_39_q_net <= pixel_bus_input_offset_0_9;
  delay_32_q_net <= pixel_bus_input_offset_0_10;
  delay_34_q_net <= pixel_bus_input_offset_0_11;
  delay_37_q_net <= pixel_bus_input_offset_0_12;
  delay_60_q_net <= pixel_bus_input_offset_1_2;
  delay_66_q_net <= pixel_bus_input_offset_1_3;
  delay_68_q_net <= pixel_bus_input_offset_1_4;
  delay_70_q_net <= pixel_bus_input_offset_1_5;
  delay_50_q_net <= pixel_bus_input_offset_1_6;
  delay_52_q_net <= pixel_bus_input_offset_1_7;
  delay_54_q_net <= pixel_bus_input_offset_1_8;
  delay_63_q_net <= pixel_bus_input_offset_1_9;
  delay_56_q_net <= pixel_bus_input_offset_1_10;
  delay_58_q_net <= pixel_bus_input_offset_1_11;
  delay_61_q_net <= pixel_bus_input_offset_1_12;
  delay_84_q_net <= pixel_bus_input_offset_2_2;
  delay_90_q_net <= pixel_bus_input_offset_2_3;
  delay_92_q_net <= pixel_bus_input_offset_2_4;
  delay_94_q_net <= pixel_bus_input_offset_2_5;
  delay_74_q_net <= pixel_bus_input_offset_2_6;
  delay_76_q_net <= pixel_bus_input_offset_2_7;
  delay_78_q_net <= pixel_bus_input_offset_2_8;
  delay_87_q_net <= pixel_bus_input_offset_2_9;
  delay_80_q_net <= pixel_bus_input_offset_2_10;
  delay_82_q_net <= pixel_bus_input_offset_2_11;
  delay_85_q_net <= pixel_bus_input_offset_2_12;
  delay_108_q_net <= pixel_bus_input_offset_3_2;
  delay_114_q_net <= pixel_bus_input_offset_3_3;
  delay_116_q_net <= pixel_bus_input_offset_3_4;
  delay_118_q_net <= pixel_bus_input_offset_3_5;
  delay_98_q_net <= pixel_bus_input_offset_3_6;
  delay_100_q_net <= pixel_bus_input_offset_3_7;
  delay_102_q_net <= pixel_bus_input_offset_3_8;
  delay_111_q_net <= pixel_bus_input_offset_3_9;
  delay_104_q_net <= pixel_bus_input_offset_3_10;
  delay_106_q_net <= pixel_bus_input_offset_3_11;
  delay_109_q_net <= pixel_bus_input_offset_3_12;
  delay_2_q_net <= pixel_bus_input_offset_4_2;
  delay_4_q_net <= pixel_bus_input_offset_4_3;
  delay_6_q_net <= pixel_bus_input_offset_4_4;
  delay_8_q_net <= pixel_bus_input_offset_4_5;
  delay_10_q_net <= pixel_bus_input_offset_4_6;
  delay_12_q_net <= pixel_bus_input_offset_4_7;
  delay_14_q_net <= pixel_bus_input_offset_4_8;
  delay_23_q_net <= pixel_bus_input_offset_4_9;
  delay_16_q_net <= pixel_bus_input_offset_4_10;
  delay_18_q_net <= pixel_bus_input_offset_4_11;
  delay_20_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_1_y_net <= valid_bus_input_5;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x0 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x0 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x0 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x0 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x0 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x0 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x0 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x0 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x0 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x0 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x0 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x1 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x1;
architecture structural of mh_accumlator_kernel_results_x1 is 
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x1 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x1;
architecture structural of mh_accumulator_offset_0_x1 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x1 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x1;
architecture structural of mh_accumulator_offset_1_x1 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x1 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x1;
architecture structural of mh_accumulator_offset_2_x1 is 
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x1 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x1;
architecture structural of mh_accumulator_offset_3_x1 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x1 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x1;
architecture structural of mh_accumulator_offset_4_x1 is 
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x1 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x1;
architecture structural of mh_multiple_and_add_offset_0_x1 is 
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x1 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x1;
architecture structural of mh_multiple_and_add_offset_1_x1 is 
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x1 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x1;
architecture structural of mh_multiple_and_add_offset_2_x1 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x1 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x1;
architecture structural of mh_multiple_and_add_offset_3_x1 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x1 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x1;
architecture structural of mh_multiple_and_add_offset_4_x1 is 
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_2 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_4 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_2;
architecture structural of mh_kernel_result_2 is 
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_48_q_net <= pixel_bus_input_offset_0_1;
  delay_72_q_net <= pixel_bus_input_offset_1_1;
  delay_96_q_net <= pixel_bus_input_offset_2_1;
  delay_0_q_net <= pixel_bus_input_offset_3_1;
  delay_22_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_0_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_60_q_net <= pixel_bus_input_offset_0_2;
  delay_66_q_net <= pixel_bus_input_offset_0_3;
  delay_68_q_net <= pixel_bus_input_offset_0_4;
  delay_70_q_net <= pixel_bus_input_offset_0_5;
  delay_50_q_net <= pixel_bus_input_offset_0_6;
  delay_52_q_net <= pixel_bus_input_offset_0_7;
  delay_54_q_net <= pixel_bus_input_offset_0_8;
  delay_63_q_net <= pixel_bus_input_offset_0_9;
  delay_56_q_net <= pixel_bus_input_offset_0_10;
  delay_58_q_net <= pixel_bus_input_offset_0_11;
  delay_61_q_net <= pixel_bus_input_offset_0_12;
  delay_84_q_net <= pixel_bus_input_offset_1_2;
  delay_90_q_net <= pixel_bus_input_offset_1_3;
  delay_92_q_net <= pixel_bus_input_offset_1_4;
  delay_94_q_net <= pixel_bus_input_offset_1_5;
  delay_74_q_net <= pixel_bus_input_offset_1_6;
  delay_76_q_net <= pixel_bus_input_offset_1_7;
  delay_78_q_net <= pixel_bus_input_offset_1_8;
  delay_87_q_net <= pixel_bus_input_offset_1_9;
  delay_80_q_net <= pixel_bus_input_offset_1_10;
  delay_82_q_net <= pixel_bus_input_offset_1_11;
  delay_85_q_net <= pixel_bus_input_offset_1_12;
  delay_108_q_net <= pixel_bus_input_offset_2_2;
  delay_114_q_net <= pixel_bus_input_offset_2_3;
  delay_116_q_net <= pixel_bus_input_offset_2_4;
  delay_118_q_net <= pixel_bus_input_offset_2_5;
  delay_98_q_net <= pixel_bus_input_offset_2_6;
  delay_100_q_net <= pixel_bus_input_offset_2_7;
  delay_102_q_net <= pixel_bus_input_offset_2_8;
  delay_111_q_net <= pixel_bus_input_offset_2_9;
  delay_104_q_net <= pixel_bus_input_offset_2_10;
  delay_106_q_net <= pixel_bus_input_offset_2_11;
  delay_109_q_net <= pixel_bus_input_offset_2_12;
  delay_2_q_net <= pixel_bus_input_offset_3_2;
  delay_4_q_net <= pixel_bus_input_offset_3_3;
  delay_6_q_net <= pixel_bus_input_offset_3_4;
  delay_8_q_net <= pixel_bus_input_offset_3_5;
  delay_10_q_net <= pixel_bus_input_offset_3_6;
  delay_12_q_net <= pixel_bus_input_offset_3_7;
  delay_14_q_net <= pixel_bus_input_offset_3_8;
  delay_23_q_net <= pixel_bus_input_offset_3_9;
  delay_16_q_net <= pixel_bus_input_offset_3_10;
  delay_18_q_net <= pixel_bus_input_offset_3_11;
  delay_20_q_net <= pixel_bus_input_offset_3_12;
  delay_36_q_net <= pixel_bus_input_offset_4_2;
  delay_42_q_net <= pixel_bus_input_offset_4_3;
  delay_44_q_net <= pixel_bus_input_offset_4_4;
  delay_46_q_net <= pixel_bus_input_offset_4_5;
  delay_26_q_net <= pixel_bus_input_offset_4_6;
  delay_28_q_net <= pixel_bus_input_offset_4_7;
  delay_30_q_net <= pixel_bus_input_offset_4_8;
  delay_39_q_net <= pixel_bus_input_offset_4_9;
  delay_32_q_net <= pixel_bus_input_offset_4_10;
  delay_34_q_net <= pixel_bus_input_offset_4_11;
  delay_37_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_1_y_net <= valid_bus_input_4;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x1 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x1 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x1 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x1 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x1 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x1 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x1 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x1 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x1 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x1 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x1 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x2 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x2;
architecture structural of mh_accumlator_kernel_results_x2 is 
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x2 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x2;
architecture structural of mh_accumulator_offset_0_x2 is 
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x2 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x2;
architecture structural of mh_accumulator_offset_1_x2 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x2 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x2;
architecture structural of mh_accumulator_offset_2_x2 is 
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x2 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x2;
architecture structural of mh_accumulator_offset_3_x2 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x2 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x2;
architecture structural of mh_accumulator_offset_4_x2 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x2 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x2;
architecture structural of mh_multiple_and_add_offset_0_x2 is 
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x2 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x2;
architecture structural of mh_multiple_and_add_offset_1_x2 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x2 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x2;
architecture structural of mh_multiple_and_add_offset_2_x2 is 
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x2 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x2;
architecture structural of mh_multiple_and_add_offset_3_x2 is 
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal ce_net : std_logic;
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x2 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x2;
architecture structural of mh_multiple_and_add_offset_4_x2 is 
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_3 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_3 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_3;
architecture structural of mh_kernel_result_3 is 
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_72_q_net <= pixel_bus_input_offset_0_1;
  delay_96_q_net <= pixel_bus_input_offset_1_1;
  delay_0_q_net <= pixel_bus_input_offset_2_1;
  delay_22_q_net <= pixel_bus_input_offset_3_1;
  delay_48_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_0_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_84_q_net <= pixel_bus_input_offset_0_2;
  delay_90_q_net <= pixel_bus_input_offset_0_3;
  delay_92_q_net <= pixel_bus_input_offset_0_4;
  delay_94_q_net <= pixel_bus_input_offset_0_5;
  delay_74_q_net <= pixel_bus_input_offset_0_6;
  delay_76_q_net <= pixel_bus_input_offset_0_7;
  delay_78_q_net <= pixel_bus_input_offset_0_8;
  delay_87_q_net <= pixel_bus_input_offset_0_9;
  delay_80_q_net <= pixel_bus_input_offset_0_10;
  delay_82_q_net <= pixel_bus_input_offset_0_11;
  delay_85_q_net <= pixel_bus_input_offset_0_12;
  delay_108_q_net <= pixel_bus_input_offset_1_2;
  delay_114_q_net <= pixel_bus_input_offset_1_3;
  delay_116_q_net <= pixel_bus_input_offset_1_4;
  delay_118_q_net <= pixel_bus_input_offset_1_5;
  delay_98_q_net <= pixel_bus_input_offset_1_6;
  delay_100_q_net <= pixel_bus_input_offset_1_7;
  delay_102_q_net <= pixel_bus_input_offset_1_8;
  delay_111_q_net <= pixel_bus_input_offset_1_9;
  delay_104_q_net <= pixel_bus_input_offset_1_10;
  delay_106_q_net <= pixel_bus_input_offset_1_11;
  delay_109_q_net <= pixel_bus_input_offset_1_12;
  delay_2_q_net <= pixel_bus_input_offset_2_2;
  delay_4_q_net <= pixel_bus_input_offset_2_3;
  delay_6_q_net <= pixel_bus_input_offset_2_4;
  delay_8_q_net <= pixel_bus_input_offset_2_5;
  delay_10_q_net <= pixel_bus_input_offset_2_6;
  delay_12_q_net <= pixel_bus_input_offset_2_7;
  delay_14_q_net <= pixel_bus_input_offset_2_8;
  delay_23_q_net <= pixel_bus_input_offset_2_9;
  delay_16_q_net <= pixel_bus_input_offset_2_10;
  delay_18_q_net <= pixel_bus_input_offset_2_11;
  delay_20_q_net <= pixel_bus_input_offset_2_12;
  delay_36_q_net <= pixel_bus_input_offset_3_2;
  delay_42_q_net <= pixel_bus_input_offset_3_3;
  delay_44_q_net <= pixel_bus_input_offset_3_4;
  delay_46_q_net <= pixel_bus_input_offset_3_5;
  delay_26_q_net <= pixel_bus_input_offset_3_6;
  delay_28_q_net <= pixel_bus_input_offset_3_7;
  delay_30_q_net <= pixel_bus_input_offset_3_8;
  delay_39_q_net <= pixel_bus_input_offset_3_9;
  delay_32_q_net <= pixel_bus_input_offset_3_10;
  delay_34_q_net <= pixel_bus_input_offset_3_11;
  delay_37_q_net <= pixel_bus_input_offset_3_12;
  delay_60_q_net <= pixel_bus_input_offset_4_2;
  delay_66_q_net <= pixel_bus_input_offset_4_3;
  delay_68_q_net <= pixel_bus_input_offset_4_4;
  delay_70_q_net <= pixel_bus_input_offset_4_5;
  delay_50_q_net <= pixel_bus_input_offset_4_6;
  delay_52_q_net <= pixel_bus_input_offset_4_7;
  delay_54_q_net <= pixel_bus_input_offset_4_8;
  delay_63_q_net <= pixel_bus_input_offset_4_9;
  delay_56_q_net <= pixel_bus_input_offset_4_10;
  delay_58_q_net <= pixel_bus_input_offset_4_11;
  delay_61_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_1_y_net <= valid_bus_input_3;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x2 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x2 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x2 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x2 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x2 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x2 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x2 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x2 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x2 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x2 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x2 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x3 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x3;
architecture structural of mh_accumlator_kernel_results_x3 is 
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x3 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x3;
architecture structural of mh_accumulator_offset_0_x3 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x3 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x3;
architecture structural of mh_accumulator_offset_1_x3 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x3 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x3;
architecture structural of mh_accumulator_offset_2_x3 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x3 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x3;
architecture structural of mh_accumulator_offset_3_x3 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x3 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x3;
architecture structural of mh_accumulator_offset_4_x3 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x3 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x3;
architecture structural of mh_multiple_and_add_offset_0_x3 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x3 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x3;
architecture structural of mh_multiple_and_add_offset_1_x3 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x3 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x3;
architecture structural of mh_multiple_and_add_offset_2_x3 is 
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x3 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x3;
architecture structural of mh_multiple_and_add_offset_3_x3 is 
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x3 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x3;
architecture structural of mh_multiple_and_add_offset_4_x3 is 
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal clk_net : std_logic;
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_4 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_2 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_4;
architecture structural of mh_kernel_result_4 is 
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_96_q_net <= pixel_bus_input_offset_0_1;
  delay_0_q_net <= pixel_bus_input_offset_1_1;
  delay_22_q_net <= pixel_bus_input_offset_2_1;
  delay_48_q_net <= pixel_bus_input_offset_3_1;
  delay_72_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_0_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_108_q_net <= pixel_bus_input_offset_0_2;
  delay_114_q_net <= pixel_bus_input_offset_0_3;
  delay_116_q_net <= pixel_bus_input_offset_0_4;
  delay_118_q_net <= pixel_bus_input_offset_0_5;
  delay_98_q_net <= pixel_bus_input_offset_0_6;
  delay_100_q_net <= pixel_bus_input_offset_0_7;
  delay_102_q_net <= pixel_bus_input_offset_0_8;
  delay_111_q_net <= pixel_bus_input_offset_0_9;
  delay_104_q_net <= pixel_bus_input_offset_0_10;
  delay_106_q_net <= pixel_bus_input_offset_0_11;
  delay_109_q_net <= pixel_bus_input_offset_0_12;
  delay_2_q_net <= pixel_bus_input_offset_1_2;
  delay_4_q_net <= pixel_bus_input_offset_1_3;
  delay_6_q_net <= pixel_bus_input_offset_1_4;
  delay_8_q_net <= pixel_bus_input_offset_1_5;
  delay_10_q_net <= pixel_bus_input_offset_1_6;
  delay_12_q_net <= pixel_bus_input_offset_1_7;
  delay_14_q_net <= pixel_bus_input_offset_1_8;
  delay_23_q_net <= pixel_bus_input_offset_1_9;
  delay_16_q_net <= pixel_bus_input_offset_1_10;
  delay_18_q_net <= pixel_bus_input_offset_1_11;
  delay_20_q_net <= pixel_bus_input_offset_1_12;
  delay_36_q_net <= pixel_bus_input_offset_2_2;
  delay_42_q_net <= pixel_bus_input_offset_2_3;
  delay_44_q_net <= pixel_bus_input_offset_2_4;
  delay_46_q_net <= pixel_bus_input_offset_2_5;
  delay_26_q_net <= pixel_bus_input_offset_2_6;
  delay_28_q_net <= pixel_bus_input_offset_2_7;
  delay_30_q_net <= pixel_bus_input_offset_2_8;
  delay_39_q_net <= pixel_bus_input_offset_2_9;
  delay_32_q_net <= pixel_bus_input_offset_2_10;
  delay_34_q_net <= pixel_bus_input_offset_2_11;
  delay_37_q_net <= pixel_bus_input_offset_2_12;
  delay_60_q_net <= pixel_bus_input_offset_3_2;
  delay_66_q_net <= pixel_bus_input_offset_3_3;
  delay_68_q_net <= pixel_bus_input_offset_3_4;
  delay_70_q_net <= pixel_bus_input_offset_3_5;
  delay_50_q_net <= pixel_bus_input_offset_3_6;
  delay_52_q_net <= pixel_bus_input_offset_3_7;
  delay_54_q_net <= pixel_bus_input_offset_3_8;
  delay_63_q_net <= pixel_bus_input_offset_3_9;
  delay_56_q_net <= pixel_bus_input_offset_3_10;
  delay_58_q_net <= pixel_bus_input_offset_3_11;
  delay_61_q_net <= pixel_bus_input_offset_3_12;
  delay_84_q_net <= pixel_bus_input_offset_4_2;
  delay_90_q_net <= pixel_bus_input_offset_4_3;
  delay_92_q_net <= pixel_bus_input_offset_4_4;
  delay_94_q_net <= pixel_bus_input_offset_4_5;
  delay_74_q_net <= pixel_bus_input_offset_4_6;
  delay_76_q_net <= pixel_bus_input_offset_4_7;
  delay_78_q_net <= pixel_bus_input_offset_4_8;
  delay_87_q_net <= pixel_bus_input_offset_4_9;
  delay_80_q_net <= pixel_bus_input_offset_4_10;
  delay_82_q_net <= pixel_bus_input_offset_4_11;
  delay_85_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_1_y_net <= valid_bus_input_2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x3 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x3 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x3 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x3 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x3 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x3 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x3 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x3 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x3 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x3 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x3 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x4 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x4;
architecture structural of mh_accumlator_kernel_results_x4 is 
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x4 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x4;
architecture structural of mh_accumulator_offset_0_x4 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x4 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x4;
architecture structural of mh_accumulator_offset_1_x4 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x4 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x4;
architecture structural of mh_accumulator_offset_2_x4 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x4 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x4;
architecture structural of mh_accumulator_offset_3_x4 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x4 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x4;
architecture structural of mh_accumulator_offset_4_x4 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x4 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x4;
architecture structural of mh_multiple_and_add_offset_0_x4 is 
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x4 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x4;
architecture structural of mh_multiple_and_add_offset_1_x4 is 
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x4 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x4;
architecture structural of mh_multiple_and_add_offset_2_x4 is 
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x4 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x4;
architecture structural of mh_multiple_and_add_offset_3_x4 is 
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x4 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x4;
architecture structural of mh_multiple_and_add_offset_4_x4 is 
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_5 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_5;
architecture structural of mh_kernel_result_5 is 
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_0_q_net <= pixel_bus_input_offset_0_1;
  delay_22_q_net <= pixel_bus_input_offset_1_1;
  delay_48_q_net <= pixel_bus_input_offset_2_1;
  delay_72_q_net <= pixel_bus_input_offset_3_1;
  delay_96_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_1_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_2_q_net <= pixel_bus_input_offset_0_2;
  delay_4_q_net <= pixel_bus_input_offset_0_3;
  delay_6_q_net <= pixel_bus_input_offset_0_4;
  delay_8_q_net <= pixel_bus_input_offset_0_5;
  delay_10_q_net <= pixel_bus_input_offset_0_6;
  delay_12_q_net <= pixel_bus_input_offset_0_7;
  delay_14_q_net <= pixel_bus_input_offset_0_8;
  delay_23_q_net <= pixel_bus_input_offset_0_9;
  delay_16_q_net <= pixel_bus_input_offset_0_10;
  delay_18_q_net <= pixel_bus_input_offset_0_11;
  delay_20_q_net <= pixel_bus_input_offset_0_12;
  delay_36_q_net <= pixel_bus_input_offset_1_2;
  delay_42_q_net <= pixel_bus_input_offset_1_3;
  delay_44_q_net <= pixel_bus_input_offset_1_4;
  delay_46_q_net <= pixel_bus_input_offset_1_5;
  delay_26_q_net <= pixel_bus_input_offset_1_6;
  delay_28_q_net <= pixel_bus_input_offset_1_7;
  delay_30_q_net <= pixel_bus_input_offset_1_8;
  delay_39_q_net <= pixel_bus_input_offset_1_9;
  delay_32_q_net <= pixel_bus_input_offset_1_10;
  delay_34_q_net <= pixel_bus_input_offset_1_11;
  delay_37_q_net <= pixel_bus_input_offset_1_12;
  delay_60_q_net <= pixel_bus_input_offset_2_2;
  delay_66_q_net <= pixel_bus_input_offset_2_3;
  delay_68_q_net <= pixel_bus_input_offset_2_4;
  delay_70_q_net <= pixel_bus_input_offset_2_5;
  delay_50_q_net <= pixel_bus_input_offset_2_6;
  delay_52_q_net <= pixel_bus_input_offset_2_7;
  delay_54_q_net <= pixel_bus_input_offset_2_8;
  delay_63_q_net <= pixel_bus_input_offset_2_9;
  delay_56_q_net <= pixel_bus_input_offset_2_10;
  delay_58_q_net <= pixel_bus_input_offset_2_11;
  delay_61_q_net <= pixel_bus_input_offset_2_12;
  delay_84_q_net <= pixel_bus_input_offset_3_2;
  delay_90_q_net <= pixel_bus_input_offset_3_3;
  delay_92_q_net <= pixel_bus_input_offset_3_4;
  delay_94_q_net <= pixel_bus_input_offset_3_5;
  delay_74_q_net <= pixel_bus_input_offset_3_6;
  delay_76_q_net <= pixel_bus_input_offset_3_7;
  delay_78_q_net <= pixel_bus_input_offset_3_8;
  delay_87_q_net <= pixel_bus_input_offset_3_9;
  delay_80_q_net <= pixel_bus_input_offset_3_10;
  delay_82_q_net <= pixel_bus_input_offset_3_11;
  delay_85_q_net <= pixel_bus_input_offset_3_12;
  delay_108_q_net <= pixel_bus_input_offset_4_2;
  delay_114_q_net <= pixel_bus_input_offset_4_3;
  delay_116_q_net <= pixel_bus_input_offset_4_4;
  delay_118_q_net <= pixel_bus_input_offset_4_5;
  delay_98_q_net <= pixel_bus_input_offset_4_6;
  delay_100_q_net <= pixel_bus_input_offset_4_7;
  delay_102_q_net <= pixel_bus_input_offset_4_8;
  delay_111_q_net <= pixel_bus_input_offset_4_9;
  delay_104_q_net <= pixel_bus_input_offset_4_10;
  delay_106_q_net <= pixel_bus_input_offset_4_11;
  delay_109_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x4 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x4 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x4 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x4 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x4 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x4 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x4 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x4 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x4 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x4 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x4 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x5 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x5;
architecture structural of mh_accumlator_kernel_results_x5 is 
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x5 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x5;
architecture structural of mh_accumulator_offset_0_x5 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x5 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x5;
architecture structural of mh_accumulator_offset_1_x5 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x5 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x5;
architecture structural of mh_accumulator_offset_2_x5 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x5 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x5;
architecture structural of mh_accumulator_offset_3_x5 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x5 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x5;
architecture structural of mh_accumulator_offset_4_x5 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x5 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x5;
architecture structural of mh_multiple_and_add_offset_0_x5 is 
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x5 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x5;
architecture structural of mh_multiple_and_add_offset_1_x5 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x5 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x5;
architecture structural of mh_multiple_and_add_offset_2_x5 is 
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x5 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x5;
architecture structural of mh_multiple_and_add_offset_3_x5 is 
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x5 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x5;
architecture structural of mh_multiple_and_add_offset_4_x5 is 
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_6 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_5 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_6;
architecture structural of mh_kernel_result_6 is 
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_22_q_net <= pixel_bus_input_offset_0_1;
  delay_48_q_net <= pixel_bus_input_offset_1_1;
  delay_72_q_net <= pixel_bus_input_offset_2_1;
  delay_96_q_net <= pixel_bus_input_offset_3_1;
  delay_0_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_1_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_36_q_net <= pixel_bus_input_offset_0_2;
  delay_42_q_net <= pixel_bus_input_offset_0_3;
  delay_44_q_net <= pixel_bus_input_offset_0_4;
  delay_46_q_net <= pixel_bus_input_offset_0_5;
  delay_26_q_net <= pixel_bus_input_offset_0_6;
  delay_28_q_net <= pixel_bus_input_offset_0_7;
  delay_30_q_net <= pixel_bus_input_offset_0_8;
  delay_39_q_net <= pixel_bus_input_offset_0_9;
  delay_32_q_net <= pixel_bus_input_offset_0_10;
  delay_34_q_net <= pixel_bus_input_offset_0_11;
  delay_37_q_net <= pixel_bus_input_offset_0_12;
  delay_60_q_net <= pixel_bus_input_offset_1_2;
  delay_66_q_net <= pixel_bus_input_offset_1_3;
  delay_68_q_net <= pixel_bus_input_offset_1_4;
  delay_70_q_net <= pixel_bus_input_offset_1_5;
  delay_50_q_net <= pixel_bus_input_offset_1_6;
  delay_52_q_net <= pixel_bus_input_offset_1_7;
  delay_54_q_net <= pixel_bus_input_offset_1_8;
  delay_63_q_net <= pixel_bus_input_offset_1_9;
  delay_56_q_net <= pixel_bus_input_offset_1_10;
  delay_58_q_net <= pixel_bus_input_offset_1_11;
  delay_61_q_net <= pixel_bus_input_offset_1_12;
  delay_84_q_net <= pixel_bus_input_offset_2_2;
  delay_90_q_net <= pixel_bus_input_offset_2_3;
  delay_92_q_net <= pixel_bus_input_offset_2_4;
  delay_94_q_net <= pixel_bus_input_offset_2_5;
  delay_74_q_net <= pixel_bus_input_offset_2_6;
  delay_76_q_net <= pixel_bus_input_offset_2_7;
  delay_78_q_net <= pixel_bus_input_offset_2_8;
  delay_87_q_net <= pixel_bus_input_offset_2_9;
  delay_80_q_net <= pixel_bus_input_offset_2_10;
  delay_82_q_net <= pixel_bus_input_offset_2_11;
  delay_85_q_net <= pixel_bus_input_offset_2_12;
  delay_108_q_net <= pixel_bus_input_offset_3_2;
  delay_114_q_net <= pixel_bus_input_offset_3_3;
  delay_116_q_net <= pixel_bus_input_offset_3_4;
  delay_118_q_net <= pixel_bus_input_offset_3_5;
  delay_98_q_net <= pixel_bus_input_offset_3_6;
  delay_100_q_net <= pixel_bus_input_offset_3_7;
  delay_102_q_net <= pixel_bus_input_offset_3_8;
  delay_111_q_net <= pixel_bus_input_offset_3_9;
  delay_104_q_net <= pixel_bus_input_offset_3_10;
  delay_106_q_net <= pixel_bus_input_offset_3_11;
  delay_109_q_net <= pixel_bus_input_offset_3_12;
  delay_2_q_net <= pixel_bus_input_offset_4_2;
  delay_4_q_net <= pixel_bus_input_offset_4_3;
  delay_6_q_net <= pixel_bus_input_offset_4_4;
  delay_8_q_net <= pixel_bus_input_offset_4_5;
  delay_10_q_net <= pixel_bus_input_offset_4_6;
  delay_12_q_net <= pixel_bus_input_offset_4_7;
  delay_14_q_net <= pixel_bus_input_offset_4_8;
  delay_23_q_net <= pixel_bus_input_offset_4_9;
  delay_16_q_net <= pixel_bus_input_offset_4_10;
  delay_18_q_net <= pixel_bus_input_offset_4_11;
  delay_20_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_0_y_net <= valid_bus_input_5;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x5 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x5 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x5 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x5 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x5 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x5 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x5 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x5 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x5 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x5 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x5 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x6 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x6;
architecture structural of mh_accumlator_kernel_results_x6 is 
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x6 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x6;
architecture structural of mh_accumulator_offset_0_x6 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x6 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x6;
architecture structural of mh_accumulator_offset_1_x6 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x6 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x6;
architecture structural of mh_accumulator_offset_2_x6 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal clk_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x6 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x6;
architecture structural of mh_accumulator_offset_3_x6 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal clk_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x6 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x6;
architecture structural of mh_accumulator_offset_4_x6 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x6 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x6;
architecture structural of mh_multiple_and_add_offset_0_x6 is 
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x6 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x6;
architecture structural of mh_multiple_and_add_offset_1_x6 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x6 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x6;
architecture structural of mh_multiple_and_add_offset_2_x6 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x6 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x6;
architecture structural of mh_multiple_and_add_offset_3_x6 is 
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x6 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x6;
architecture structural of mh_multiple_and_add_offset_4_x6 is 
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_7 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_4 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_7;
architecture structural of mh_kernel_result_7 is 
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_48_q_net <= pixel_bus_input_offset_0_1;
  delay_72_q_net <= pixel_bus_input_offset_1_1;
  delay_96_q_net <= pixel_bus_input_offset_2_1;
  delay_0_q_net <= pixel_bus_input_offset_3_1;
  delay_22_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_1_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_60_q_net <= pixel_bus_input_offset_0_2;
  delay_66_q_net <= pixel_bus_input_offset_0_3;
  delay_68_q_net <= pixel_bus_input_offset_0_4;
  delay_70_q_net <= pixel_bus_input_offset_0_5;
  delay_50_q_net <= pixel_bus_input_offset_0_6;
  delay_52_q_net <= pixel_bus_input_offset_0_7;
  delay_54_q_net <= pixel_bus_input_offset_0_8;
  delay_63_q_net <= pixel_bus_input_offset_0_9;
  delay_56_q_net <= pixel_bus_input_offset_0_10;
  delay_58_q_net <= pixel_bus_input_offset_0_11;
  delay_61_q_net <= pixel_bus_input_offset_0_12;
  delay_84_q_net <= pixel_bus_input_offset_1_2;
  delay_90_q_net <= pixel_bus_input_offset_1_3;
  delay_92_q_net <= pixel_bus_input_offset_1_4;
  delay_94_q_net <= pixel_bus_input_offset_1_5;
  delay_74_q_net <= pixel_bus_input_offset_1_6;
  delay_76_q_net <= pixel_bus_input_offset_1_7;
  delay_78_q_net <= pixel_bus_input_offset_1_8;
  delay_87_q_net <= pixel_bus_input_offset_1_9;
  delay_80_q_net <= pixel_bus_input_offset_1_10;
  delay_82_q_net <= pixel_bus_input_offset_1_11;
  delay_85_q_net <= pixel_bus_input_offset_1_12;
  delay_108_q_net <= pixel_bus_input_offset_2_2;
  delay_114_q_net <= pixel_bus_input_offset_2_3;
  delay_116_q_net <= pixel_bus_input_offset_2_4;
  delay_118_q_net <= pixel_bus_input_offset_2_5;
  delay_98_q_net <= pixel_bus_input_offset_2_6;
  delay_100_q_net <= pixel_bus_input_offset_2_7;
  delay_102_q_net <= pixel_bus_input_offset_2_8;
  delay_111_q_net <= pixel_bus_input_offset_2_9;
  delay_104_q_net <= pixel_bus_input_offset_2_10;
  delay_106_q_net <= pixel_bus_input_offset_2_11;
  delay_109_q_net <= pixel_bus_input_offset_2_12;
  delay_2_q_net <= pixel_bus_input_offset_3_2;
  delay_4_q_net <= pixel_bus_input_offset_3_3;
  delay_6_q_net <= pixel_bus_input_offset_3_4;
  delay_8_q_net <= pixel_bus_input_offset_3_5;
  delay_10_q_net <= pixel_bus_input_offset_3_6;
  delay_12_q_net <= pixel_bus_input_offset_3_7;
  delay_14_q_net <= pixel_bus_input_offset_3_8;
  delay_23_q_net <= pixel_bus_input_offset_3_9;
  delay_16_q_net <= pixel_bus_input_offset_3_10;
  delay_18_q_net <= pixel_bus_input_offset_3_11;
  delay_20_q_net <= pixel_bus_input_offset_3_12;
  delay_36_q_net <= pixel_bus_input_offset_4_2;
  delay_42_q_net <= pixel_bus_input_offset_4_3;
  delay_44_q_net <= pixel_bus_input_offset_4_4;
  delay_46_q_net <= pixel_bus_input_offset_4_5;
  delay_26_q_net <= pixel_bus_input_offset_4_6;
  delay_28_q_net <= pixel_bus_input_offset_4_7;
  delay_30_q_net <= pixel_bus_input_offset_4_8;
  delay_39_q_net <= pixel_bus_input_offset_4_9;
  delay_32_q_net <= pixel_bus_input_offset_4_10;
  delay_34_q_net <= pixel_bus_input_offset_4_11;
  delay_37_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_0_y_net <= valid_bus_input_4;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x6 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x6 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x6 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x6 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x6 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x6 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x6 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x6 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x6 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x6 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x6 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x7 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x7;
architecture structural of mh_accumlator_kernel_results_x7 is 
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x7 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x7;
architecture structural of mh_accumulator_offset_0_x7 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x7 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x7;
architecture structural of mh_accumulator_offset_1_x7 is 
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x7 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x7;
architecture structural of mh_accumulator_offset_2_x7 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal ce_net : std_logic;
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x7 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x7;
architecture structural of mh_accumulator_offset_3_x7 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x7 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x7;
architecture structural of mh_accumulator_offset_4_x7 is 
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x7 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x7;
architecture structural of mh_multiple_and_add_offset_0_x7 is 
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x7 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x7;
architecture structural of mh_multiple_and_add_offset_1_x7 is 
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x7 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x7;
architecture structural of mh_multiple_and_add_offset_2_x7 is 
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal ce_net : std_logic;
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x7 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x7;
architecture structural of mh_multiple_and_add_offset_3_x7 is 
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x7 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x7;
architecture structural of mh_multiple_and_add_offset_4_x7 is 
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal clk_net : std_logic;
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 8
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_8 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_3 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_8;
architecture structural of mh_kernel_result_8 is 
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_72_q_net <= pixel_bus_input_offset_0_1;
  delay_96_q_net <= pixel_bus_input_offset_1_1;
  delay_0_q_net <= pixel_bus_input_offset_2_1;
  delay_22_q_net <= pixel_bus_input_offset_3_1;
  delay_48_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_1_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_84_q_net <= pixel_bus_input_offset_0_2;
  delay_90_q_net <= pixel_bus_input_offset_0_3;
  delay_92_q_net <= pixel_bus_input_offset_0_4;
  delay_94_q_net <= pixel_bus_input_offset_0_5;
  delay_74_q_net <= pixel_bus_input_offset_0_6;
  delay_76_q_net <= pixel_bus_input_offset_0_7;
  delay_78_q_net <= pixel_bus_input_offset_0_8;
  delay_87_q_net <= pixel_bus_input_offset_0_9;
  delay_80_q_net <= pixel_bus_input_offset_0_10;
  delay_82_q_net <= pixel_bus_input_offset_0_11;
  delay_85_q_net <= pixel_bus_input_offset_0_12;
  delay_108_q_net <= pixel_bus_input_offset_1_2;
  delay_114_q_net <= pixel_bus_input_offset_1_3;
  delay_116_q_net <= pixel_bus_input_offset_1_4;
  delay_118_q_net <= pixel_bus_input_offset_1_5;
  delay_98_q_net <= pixel_bus_input_offset_1_6;
  delay_100_q_net <= pixel_bus_input_offset_1_7;
  delay_102_q_net <= pixel_bus_input_offset_1_8;
  delay_111_q_net <= pixel_bus_input_offset_1_9;
  delay_104_q_net <= pixel_bus_input_offset_1_10;
  delay_106_q_net <= pixel_bus_input_offset_1_11;
  delay_109_q_net <= pixel_bus_input_offset_1_12;
  delay_2_q_net <= pixel_bus_input_offset_2_2;
  delay_4_q_net <= pixel_bus_input_offset_2_3;
  delay_6_q_net <= pixel_bus_input_offset_2_4;
  delay_8_q_net <= pixel_bus_input_offset_2_5;
  delay_10_q_net <= pixel_bus_input_offset_2_6;
  delay_12_q_net <= pixel_bus_input_offset_2_7;
  delay_14_q_net <= pixel_bus_input_offset_2_8;
  delay_23_q_net <= pixel_bus_input_offset_2_9;
  delay_16_q_net <= pixel_bus_input_offset_2_10;
  delay_18_q_net <= pixel_bus_input_offset_2_11;
  delay_20_q_net <= pixel_bus_input_offset_2_12;
  delay_36_q_net <= pixel_bus_input_offset_3_2;
  delay_42_q_net <= pixel_bus_input_offset_3_3;
  delay_44_q_net <= pixel_bus_input_offset_3_4;
  delay_46_q_net <= pixel_bus_input_offset_3_5;
  delay_26_q_net <= pixel_bus_input_offset_3_6;
  delay_28_q_net <= pixel_bus_input_offset_3_7;
  delay_30_q_net <= pixel_bus_input_offset_3_8;
  delay_39_q_net <= pixel_bus_input_offset_3_9;
  delay_32_q_net <= pixel_bus_input_offset_3_10;
  delay_34_q_net <= pixel_bus_input_offset_3_11;
  delay_37_q_net <= pixel_bus_input_offset_3_12;
  delay_60_q_net <= pixel_bus_input_offset_4_2;
  delay_66_q_net <= pixel_bus_input_offset_4_3;
  delay_68_q_net <= pixel_bus_input_offset_4_4;
  delay_70_q_net <= pixel_bus_input_offset_4_5;
  delay_50_q_net <= pixel_bus_input_offset_4_6;
  delay_52_q_net <= pixel_bus_input_offset_4_7;
  delay_54_q_net <= pixel_bus_input_offset_4_8;
  delay_63_q_net <= pixel_bus_input_offset_4_9;
  delay_56_q_net <= pixel_bus_input_offset_4_10;
  delay_58_q_net <= pixel_bus_input_offset_4_11;
  delay_61_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_0_y_net <= valid_bus_input_3;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x7 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x7 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x7 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x7 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x7 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x7 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x7 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x7 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x7 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x7 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x7 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Accumlator Kernel Results
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumlator_kernel_results_x8 is
  port (
    slice_input_0 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_0 : in std_logic_vector( 1-1 downto 0 );
    slice_input_1 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_1 : in std_logic_vector( 1-1 downto 0 );
    slice_input_2 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_2 : in std_logic_vector( 1-1 downto 0 );
    slice_input_3 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_3 : in std_logic_vector( 1-1 downto 0 );
    slice_input_4 : in std_logic_vector( 64-1 downto 0 );
    slice_enable_4 : in std_logic_vector( 1-1 downto 0 );
    reset_collector : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumlator_kernel_results_x8;
architecture structural of mh_accumlator_kernel_results_x8 is 
  signal enable_up1_y_net : std_logic_vector( 1-1 downto 0 );
  signal result_is_valid_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_1_s_net : std_logic_vector( 65-1 downto 0 );
  signal enable_or_slice_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 64-1 downto 0 );
  signal added_slice_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 64-1 downto 0 );
  signal addition_2_s_net : std_logic_vector( 66-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 64-1 downto 0 );
  signal enable_or_slice_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal added_slice_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_or_slice_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addition_0_s_net : std_logic_vector( 65-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 64-1 downto 0 );
  signal added_slice_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 64-1 downto 0 );
  signal convert_to_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 64-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
  signal delay_enable_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_up_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_enable_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal addition_3_s_net : std_logic_vector( 67-1 downto 0 );
  signal hard_reset_y_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_3_q_net : std_logic_vector( 67-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  accumulator_0_q_net <= slice_input_0;
  delay2_q_net <= slice_enable_0;
  accumulator_0_q_net_x0 <= slice_input_1;
  delay2_q_net_x0 <= slice_enable_1;
  accumulator_0_q_net_x1 <= slice_input_2;
  delay2_q_net_x1 <= slice_enable_2;
  accumulator_0_q_net_x2 <= slice_input_3;
  delay2_q_net_x2 <= slice_enable_3;
  accumulator_0_q_net_x3 <= slice_input_4;
  delay2_q_net_x3 <= slice_enable_4;
  delay_addition8_q_net <= reset_collector;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_kernel_result_0 : entity xil_defaultlib.sysgen_accum_6061dd473e 
  port map (
    clr => '0',
    b => delay_enable_3_q_net,
    rst => hard_reset_y_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_kernel_result_0_q_net
  );
  added_slice_0 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_0_op_net
  );
  added_slice_1 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_1_op_net
  );
  added_slice_2 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_2_op_net
  );
  added_slice_3 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_3_op_net
  );
  added_slice_4 : entity xil_defaultlib.sysgen_counter_80cc42ed60 
  port map (
    clr => '0',
    en => enable_or_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => added_slice_4_op_net
  );
  addition_0 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_0_y_net,
    b => mux_slice_1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_0_s_net
  );
  addition_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 64,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 65,
    core_name0 => "mh_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 65,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 65
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_slice_2_y_net,
    b => mux_slice_3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_1_s_net
  );
  addition_2 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 65,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 65,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 66,
    core_name0 => "mh_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 66,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 66
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_0_s_net,
    b => addition_1_s_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_2_s_net
  );
  addition_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 66,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 64,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 67,
    core_name0 => "mh_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 67,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 67
  )
  port map (
    clr => '0',
    en => "1",
    a => addition_2_s_net,
    b => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addition_3_s_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  convert_to_bool_0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_0_op_net,
    y => convert_to_bool_0_y_net
  );
  convert_to_bool_1 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_1_op_net,
    y => convert_to_bool_1_y_net
  );
  convert_to_bool_2 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_2_op_net,
    y => convert_to_bool_2_y_net
  );
  convert_to_bool_3 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_3_op_net,
    y => convert_to_bool_3_y_net
  );
  convert_to_bool_4 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 1,
    y_width => 1
  )
  port map (
    x => added_slice_4_op_net,
    y => convert_to_bool_4_y_net
  );
  delay_addition_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_slice_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_0_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 64
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_enable_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_up_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_0_q_net
  );
  delay_enable_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_1_q_net
  );
  delay_enable_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_2_q_net
  );
  delay_enable_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 67
  )
  port map (
    en => '1',
    rst => '0',
    d => addition_3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_3_q_net
  );
  delay_enable_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_enable_4_q_net
  );
  enable_or_slice_0 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_0_y_net
  );
  enable_or_slice_1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x0,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_1_y_net
  );
  enable_or_slice_2 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x1,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_2_y_net
  );
  enable_or_slice_3 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x2,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_3_y_net
  );
  enable_or_slice_4 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay2_q_net_x3,
    d1 => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_or_slice_4_y_net
  );
  enable_up : entity xil_defaultlib.sysgen_logical_dcdc89c7c2 
  port map (
    clr => '0',
    d0 => delay2_q_net,
    d1 => delay2_q_net_x0,
    d2 => delay2_q_net_x1,
    d3 => delay2_q_net_x2,
    d4 => delay2_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => enable_up_y_net
  );
  enable_up1 : entity xil_defaultlib.sysgen_logical_214b4eae2b 
  port map (
    clr => '0',
    d0 => convert_to_bool_0_y_net,
    d1 => convert_to_bool_1_y_net,
    d2 => convert_to_bool_2_y_net,
    d3 => convert_to_bool_3_y_net,
    d4 => convert_to_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_up1_y_net
  );
  hard_reset : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => result_is_valid_y_net,
    clk => clk_net,
    ce => ce_net,
    y => hard_reset_y_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_bdbe110a88 
  port map (
    clr => '0',
    sel => delay2_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  result_is_valid : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_enable_2_q_net,
    d1 => enable_up1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => result_is_valid_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Accumulator Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_0_x8 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_0_x8;
architecture structural of mh_accumulator_offset_0_x8 is 
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Accumulator Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_1_x8 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_1_x8;
architecture structural of mh_accumulator_offset_1_x8 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Accumulator Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_2_x8 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_2_x8;
architecture structural of mh_accumulator_offset_2_x8 is 
  signal ce_net : std_logic;
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Accumulator Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_3_x8 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_3_x8;
architecture structural of mh_accumulator_offset_3_x8 is 
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Accumulator Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_accumulator_offset_4_x8 is
  port (
    input_value : in std_logic_vector( 34-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    last_row : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    accumulator_output : out std_logic_vector( 64-1 downto 0 );
    accumulator_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_accumulator_offset_4_x8;
architecture structural of mh_accumulator_offset_4_x8 is 
  signal ce_net : std_logic;
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  accumulator_output <= accumulator_0_q_net;
  accumulator_valid <= delay2_q_net;
  last_combine_s_net <= input_value;
  delay_addition4_q_net <= input_valid;
  delay_addition4_q_net_x0 <= last_row;
  delay_addition8_q_net <= hard_reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumulator_0 : entity xil_defaultlib.sysgen_accum_2292eb0fee 
  port map (
    clr => '0',
    b => mux_y_net,
    rst => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_0_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_8eb6000ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay_addition4_q_net,
    d1 => delay_addition4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => delay_addition8_q_net,
    d1 => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  mux : entity xil_defaultlib.sysgen_mux_d82735c294 
  port map (
    clr => '0',
    sel => delay_addition4_q_net,
    d0 => constant_op_net,
    d1 => last_combine_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Multiple and Add Offset 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_0_x8 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_0_x8;
architecture structural of mh_multiple_and_add_offset_0_x8 is 
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_96_q_net <= pixel_0;
  delay_1_q_net <= weight_0;
  delay_108_q_net <= pixel_1;
  delay_3_q_net <= weight_1;
  delay_114_q_net <= pixel_2;
  delay_5_q_net <= weight_2;
  delay_116_q_net <= pixel_3;
  delay_7_q_net <= weight_3;
  delay_118_q_net <= pixel_4;
  delay_9_q_net <= weight_4;
  delay_98_q_net <= pixel_5;
  delay_11_q_net <= weight_5;
  delay_100_q_net <= pixel_6;
  delay_13_q_net <= weight_6;
  delay_102_q_net <= pixel_7;
  delay_15_q_net <= weight_7;
  delay_111_q_net <= pixel_8;
  delay_24_q_net <= weight_8;
  delay_104_q_net <= pixel_9;
  delay_17_q_net <= weight_9;
  delay_106_q_net <= pixel_10;
  delay_19_q_net <= weight_10;
  delay_109_q_net <= pixel_11;
  delay_21_q_net <= weight_11;
  enable_passthrough_case_1_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_96_q_net,
    b => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_108_q_net,
    b => delay_3_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_106_q_net,
    b => delay_19_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_109_q_net,
    b => delay_21_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_114_q_net,
    b => delay_5_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_116_q_net,
    b => delay_7_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_118_q_net,
    b => delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_98_q_net,
    b => delay_11_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_100_q_net,
    b => delay_13_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_102_q_net,
    b => delay_15_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_111_q_net,
    b => delay_24_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_104_q_net,
    b => delay_17_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Multiple and Add Offset 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_1_x8 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_1_x8;
architecture structural of mh_multiple_and_add_offset_1_x8 is 
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_0_q_net <= pixel_0;
  delay_25_q_net <= weight_0;
  delay_2_q_net <= pixel_1;
  delay_41_q_net <= weight_1;
  delay_4_q_net <= pixel_2;
  delay_43_q_net <= weight_2;
  delay_6_q_net <= pixel_3;
  delay_45_q_net <= weight_3;
  delay_8_q_net <= pixel_4;
  delay_47_q_net <= weight_4;
  delay_10_q_net <= pixel_5;
  delay_27_q_net <= weight_5;
  delay_12_q_net <= pixel_6;
  delay_29_q_net <= weight_6;
  delay_14_q_net <= pixel_7;
  delay_31_q_net <= weight_7;
  delay_23_q_net <= pixel_8;
  delay_40_q_net <= weight_8;
  delay_16_q_net <= pixel_9;
  delay_33_q_net <= weight_9;
  delay_18_q_net <= pixel_10;
  delay_35_q_net <= weight_10;
  delay_20_q_net <= pixel_11;
  delay_38_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_0_q_net,
    b => delay_25_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_2_q_net,
    b => delay_41_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_18_q_net,
    b => delay_35_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_20_q_net,
    b => delay_38_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_4_q_net,
    b => delay_43_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_6_q_net,
    b => delay_45_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_8_q_net,
    b => delay_47_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_10_q_net,
    b => delay_27_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_12_q_net,
    b => delay_29_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_14_q_net,
    b => delay_31_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_23_q_net,
    b => delay_40_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_16_q_net,
    b => delay_33_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Multiple and Add Offset 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_2_x8 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_2_x8;
architecture structural of mh_multiple_and_add_offset_2_x8 is 
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_22_q_net <= pixel_0;
  delay_49_q_net <= weight_0;
  delay_36_q_net <= pixel_1;
  delay_65_q_net <= weight_1;
  delay_42_q_net <= pixel_2;
  delay_67_q_net <= weight_2;
  delay_44_q_net <= pixel_3;
  delay_69_q_net <= weight_3;
  delay_46_q_net <= pixel_4;
  delay_71_q_net <= weight_4;
  delay_26_q_net <= pixel_5;
  delay_51_q_net <= weight_5;
  delay_28_q_net <= pixel_6;
  delay_53_q_net <= weight_6;
  delay_30_q_net <= pixel_7;
  delay_55_q_net <= weight_7;
  delay_39_q_net <= pixel_8;
  delay_64_q_net <= weight_8;
  delay_32_q_net <= pixel_9;
  delay_57_q_net <= weight_9;
  delay_34_q_net <= pixel_10;
  delay_59_q_net <= weight_10;
  delay_37_q_net <= pixel_11;
  delay_62_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_22_q_net,
    b => delay_49_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_36_q_net,
    b => delay_65_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_34_q_net,
    b => delay_59_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_37_q_net,
    b => delay_62_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_42_q_net,
    b => delay_67_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_44_q_net,
    b => delay_69_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_46_q_net,
    b => delay_71_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_26_q_net,
    b => delay_51_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_28_q_net,
    b => delay_53_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_30_q_net,
    b => delay_55_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_39_q_net,
    b => delay_64_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_32_q_net,
    b => delay_57_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Multiple and Add Offset 3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_3_x8 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_3_x8;
architecture structural of mh_multiple_and_add_offset_3_x8 is 
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_48_q_net <= pixel_0;
  delay_73_q_net <= weight_0;
  delay_60_q_net <= pixel_1;
  delay_89_q_net <= weight_1;
  delay_66_q_net <= pixel_2;
  delay_91_q_net <= weight_2;
  delay_68_q_net <= pixel_3;
  delay_93_q_net <= weight_3;
  delay_70_q_net <= pixel_4;
  delay_95_q_net <= weight_4;
  delay_50_q_net <= pixel_5;
  delay_75_q_net <= weight_5;
  delay_52_q_net <= pixel_6;
  delay_77_q_net <= weight_6;
  delay_54_q_net <= pixel_7;
  delay_79_q_net <= weight_7;
  delay_63_q_net <= pixel_8;
  delay_88_q_net <= weight_8;
  delay_56_q_net <= pixel_9;
  delay_81_q_net <= weight_9;
  delay_58_q_net <= pixel_10;
  delay_83_q_net <= weight_10;
  delay_61_q_net <= pixel_11;
  delay_86_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_48_q_net,
    b => delay_73_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_60_q_net,
    b => delay_89_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_58_q_net,
    b => delay_83_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_61_q_net,
    b => delay_86_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_66_q_net,
    b => delay_91_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_68_q_net,
    b => delay_93_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_70_q_net,
    b => delay_95_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_50_q_net,
    b => delay_75_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_52_q_net,
    b => delay_77_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_54_q_net,
    b => delay_79_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_63_q_net,
    b => delay_88_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_56_q_net,
    b => delay_81_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9/Multiple and Add Offset 4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_multiple_and_add_offset_4_x8 is
  port (
    pixel_0 : in std_logic_vector( 12-1 downto 0 );
    weight_0 : in std_logic_vector( 18-1 downto 0 );
    pixel_1 : in std_logic_vector( 12-1 downto 0 );
    weight_1 : in std_logic_vector( 18-1 downto 0 );
    pixel_2 : in std_logic_vector( 12-1 downto 0 );
    weight_2 : in std_logic_vector( 18-1 downto 0 );
    pixel_3 : in std_logic_vector( 12-1 downto 0 );
    weight_3 : in std_logic_vector( 18-1 downto 0 );
    pixel_4 : in std_logic_vector( 12-1 downto 0 );
    weight_4 : in std_logic_vector( 18-1 downto 0 );
    pixel_5 : in std_logic_vector( 12-1 downto 0 );
    weight_5 : in std_logic_vector( 18-1 downto 0 );
    pixel_6 : in std_logic_vector( 12-1 downto 0 );
    weight_6 : in std_logic_vector( 18-1 downto 0 );
    pixel_7 : in std_logic_vector( 12-1 downto 0 );
    weight_7 : in std_logic_vector( 18-1 downto 0 );
    pixel_8 : in std_logic_vector( 12-1 downto 0 );
    weight_8 : in std_logic_vector( 18-1 downto 0 );
    pixel_9 : in std_logic_vector( 12-1 downto 0 );
    weight_9 : in std_logic_vector( 18-1 downto 0 );
    pixel_10 : in std_logic_vector( 12-1 downto 0 );
    weight_10 : in std_logic_vector( 18-1 downto 0 );
    pixel_11 : in std_logic_vector( 12-1 downto 0 );
    weight_11 : in std_logic_vector( 18-1 downto 0 );
    valid_data : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    slice_out : out std_logic_vector( 34-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end mh_multiple_and_add_offset_4_x8;
architecture structural of mh_multiple_and_add_offset_4_x8 is 
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_8_9_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_10_11_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_4_5_6_7_s_net : std_logic_vector( 33-1 downto 0 );
  signal combine_2_3_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal combine_0_1_s_net : std_logic_vector( 31-1 downto 0 );
  signal combine_0_1_2_3_s_net : std_logic_vector( 32-1 downto 0 );
  signal combine_6_7_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal pixel_0_x_weight_0_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_1_x_weight_1_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal combine_4_5_s_net : std_logic_vector( 31-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal combine_8_9_10_11_s_net : std_logic_vector( 32-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal combine_4_5_6_7_s_net : std_logic_vector( 32-1 downto 0 );
  signal pixel_10_x_weight_10_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_q_net : std_logic_vector( 32-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal pixel_11_x_weight_11_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_2_x_weight_2_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_4_x_weight_4_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_7_x_weight_7_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_3_x_weight_3_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_5_x_weight_5_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_6_x_weight_6_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_9_x_weight_9_p_net : std_logic_vector( 30-1 downto 0 );
  signal pixel_8_x_weight_8_p_net : std_logic_vector( 30-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  slice_out <= last_combine_s_net;
  valid_out <= delay_addition4_q_net;
  delay_72_q_net <= pixel_0;
  delay_97_q_net <= weight_0;
  delay_84_q_net <= pixel_1;
  delay_113_q_net <= weight_1;
  delay_90_q_net <= pixel_2;
  delay_115_q_net <= weight_2;
  delay_92_q_net <= pixel_3;
  delay_117_q_net <= weight_3;
  delay_94_q_net <= pixel_4;
  delay_119_q_net <= weight_4;
  delay_74_q_net <= pixel_5;
  delay_99_q_net <= weight_5;
  delay_76_q_net <= pixel_6;
  delay_101_q_net <= weight_6;
  delay_78_q_net <= pixel_7;
  delay_103_q_net <= weight_7;
  delay_87_q_net <= pixel_8;
  delay_112_q_net <= weight_8;
  delay_80_q_net <= pixel_9;
  delay_105_q_net <= weight_9;
  delay_82_q_net <= pixel_10;
  delay_107_q_net <= weight_10;
  delay_85_q_net <= pixel_11;
  delay_110_q_net <= weight_11;
  enable_passthrough_case_0_y_net <= valid_data;
  clk_net <= clk_1;
  ce_net <= ce_1;
  combine_0_1_2_3_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 32,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 33,
    core_name0 => "mh_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 33,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 33
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_s_net,
    b => combine_4_5_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_4_5_6_7_s_net
  );
  combine_0_1_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_s_net,
    b => combine_2_3_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_2_3_s_net
  );
  combine_4_5_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_4_5_s_net,
    b => combine_6_7_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_6_7_s_net
  );
  combine_8_9_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 31,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 31,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 32,
    core_name0 => "mh_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 32,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 32
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_8_9_s_net,
    b => combine_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_10_11_s_net
  );
  combine_0_1 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_0_x_weight_0_p_net,
    b => pixel_1_x_weight_1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_0_1_s_net
  );
  combine_10_11 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_10_x_weight_10_p_net,
    b => pixel_11_x_weight_11_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_10_11_s_net
  );
  combine_2_3 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_2_x_weight_2_p_net,
    b => pixel_3_x_weight_3_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_2_3_s_net
  );
  combine_4_5 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_4_x_weight_4_p_net,
    b => pixel_5_x_weight_5_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_4_5_s_net
  );
  combine_6_7 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_6_x_weight_6_p_net,
    b => pixel_7_x_weight_7_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_6_7_s_net
  );
  combine_8_9 : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 30,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 30,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 31,
    core_name0 => "mh_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 31,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 31
  )
  port map (
    clr => '0',
    en => "1",
    a => pixel_8_x_weight_8_p_net,
    b => pixel_9_x_weight_9_p_net,
    clk => clk_net,
    ce => ce_net,
    s => combine_8_9_s_net
  );
  delay_addition : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 32
  )
  port map (
    en => '1',
    rst => '0',
    d => combine_8_9_10_11_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_passthrough_case_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net
  );
  last_combine : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 33,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 32,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 34,
    core_name0 => "mh_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 34,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 34
  )
  port map (
    clr => '0',
    en => "1",
    a => combine_0_1_2_3_4_5_6_7_s_net,
    b => delay_addition_q_net,
    clk => clk_net,
    ce => ce_net,
    s => last_combine_s_net
  );
  pixel_0_x_weight_0 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_72_q_net,
    b => delay_97_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_0_x_weight_0_p_net
  );
  pixel_1_x_weight_1 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_84_q_net,
    b => delay_113_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_1_x_weight_1_p_net
  );
  pixel_10_x_weight_10 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_82_q_net,
    b => delay_107_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_10_x_weight_10_p_net
  );
  pixel_11_x_weight_11 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_85_q_net,
    b => delay_110_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_11_x_weight_11_p_net
  );
  pixel_2_x_weight_2 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_90_q_net,
    b => delay_115_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_2_x_weight_2_p_net
  );
  pixel_3_x_weight_3 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_92_q_net,
    b => delay_117_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_3_x_weight_3_p_net
  );
  pixel_4_x_weight_4 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_94_q_net,
    b => delay_119_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_4_x_weight_4_p_net
  );
  pixel_5_x_weight_5 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_74_q_net,
    b => delay_99_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_5_x_weight_5_p_net
  );
  pixel_6_x_weight_6 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_76_q_net,
    b => delay_101_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_6_x_weight_6_p_net
  );
  pixel_7_x_weight_7 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_78_q_net,
    b => delay_103_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_7_x_weight_7_p_net
  );
  pixel_8_x_weight_8 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_87_q_net,
    b => delay_112_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_8_x_weight_8_p_net
  );
  pixel_9_x_weight_9 : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 12,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_a_type => 1,
    c_a_width => 12,
    c_b_type => 1,
    c_b_width => 18,
    c_baat => 12,
    c_output_width => 30,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 30,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_80_q_net,
    b => delay_105_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => pixel_9_x_weight_9_p_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Kernel Result 9
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_result_9 is
  port (
    pixel_bus_input_offset_0_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_1 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_1 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_1 : in std_logic_vector( 18-1 downto 0 );
    valid_bus_input_1 : in std_logic_vector( 1-1 downto 0 );
    hard_reset : in std_logic_vector( 1-1 downto 0 );
    pixel_bus_input_offset_0_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_0_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_1_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_2_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_3_12 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_2 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_3 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_4 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_5 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_6 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_7 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_8 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_9 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_10 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_11 : in std_logic_vector( 12-1 downto 0 );
    pixel_bus_input_offset_4_12 : in std_logic_vector( 12-1 downto 0 );
    weight_bus_input_2 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_3 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_4 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_5 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_6 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_7 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_8 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_9 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_10 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_11 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_12 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_13 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_14 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_15 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_16 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_17 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_18 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_19 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_20 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_21 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_22 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_23 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_24 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_25 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_26 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_27 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_28 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_29 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_30 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_31 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_32 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_33 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_34 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_35 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_36 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_37 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_38 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_39 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_40 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_41 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_42 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_43 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_44 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_45 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_46 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_47 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_48 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_49 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_50 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_51 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_52 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_53 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_54 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_55 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_56 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_57 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_58 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_59 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_60 : in std_logic_vector( 18-1 downto 0 );
    weight_bus_input_61 : in std_logic_vector( 1-1 downto 0 );
    valid_bus_input_2 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_result_9;
architecture structural of mh_kernel_result_9 is 
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition5_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_combine_s_net_x3 : std_logic_vector( 34-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x2 : std_logic_vector( 64-1 downto 0 );
  signal accumulator_0_q_net_x0 : std_logic_vector( 64-1 downto 0 );
  signal last_combine_s_net_x1 : std_logic_vector( 34-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net_x3 : std_logic_vector( 64-1 downto 0 );
  signal delay2_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x0 : std_logic_vector( 34-1 downto 0 );
  signal last_combine_s_net : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_0_q_net_x1 : std_logic_vector( 64-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_0_q_net : std_logic_vector( 64-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal last_combine_s_net_x2 : std_logic_vector( 34-1 downto 0 );
  signal delay_addition4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay_addition4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_addition1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_addition6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= accumulator_kernel_result_0_q_net;
  valid_kernel_output <= delay_enable_4_q_net;
  delay_96_q_net <= pixel_bus_input_offset_0_1;
  delay_0_q_net <= pixel_bus_input_offset_1_1;
  delay_22_q_net <= pixel_bus_input_offset_2_1;
  delay_48_q_net <= pixel_bus_input_offset_3_1;
  delay_72_q_net <= pixel_bus_input_offset_4_1;
  delay_1_q_net <= weight_bus_input_1;
  enable_passthrough_case_1_y_net <= valid_bus_input_1;
  switch_to_zero_y_net <= hard_reset;
  delay_108_q_net <= pixel_bus_input_offset_0_2;
  delay_114_q_net <= pixel_bus_input_offset_0_3;
  delay_116_q_net <= pixel_bus_input_offset_0_4;
  delay_118_q_net <= pixel_bus_input_offset_0_5;
  delay_98_q_net <= pixel_bus_input_offset_0_6;
  delay_100_q_net <= pixel_bus_input_offset_0_7;
  delay_102_q_net <= pixel_bus_input_offset_0_8;
  delay_111_q_net <= pixel_bus_input_offset_0_9;
  delay_104_q_net <= pixel_bus_input_offset_0_10;
  delay_106_q_net <= pixel_bus_input_offset_0_11;
  delay_109_q_net <= pixel_bus_input_offset_0_12;
  delay_2_q_net <= pixel_bus_input_offset_1_2;
  delay_4_q_net <= pixel_bus_input_offset_1_3;
  delay_6_q_net <= pixel_bus_input_offset_1_4;
  delay_8_q_net <= pixel_bus_input_offset_1_5;
  delay_10_q_net <= pixel_bus_input_offset_1_6;
  delay_12_q_net <= pixel_bus_input_offset_1_7;
  delay_14_q_net <= pixel_bus_input_offset_1_8;
  delay_23_q_net <= pixel_bus_input_offset_1_9;
  delay_16_q_net <= pixel_bus_input_offset_1_10;
  delay_18_q_net <= pixel_bus_input_offset_1_11;
  delay_20_q_net <= pixel_bus_input_offset_1_12;
  delay_36_q_net <= pixel_bus_input_offset_2_2;
  delay_42_q_net <= pixel_bus_input_offset_2_3;
  delay_44_q_net <= pixel_bus_input_offset_2_4;
  delay_46_q_net <= pixel_bus_input_offset_2_5;
  delay_26_q_net <= pixel_bus_input_offset_2_6;
  delay_28_q_net <= pixel_bus_input_offset_2_7;
  delay_30_q_net <= pixel_bus_input_offset_2_8;
  delay_39_q_net <= pixel_bus_input_offset_2_9;
  delay_32_q_net <= pixel_bus_input_offset_2_10;
  delay_34_q_net <= pixel_bus_input_offset_2_11;
  delay_37_q_net <= pixel_bus_input_offset_2_12;
  delay_60_q_net <= pixel_bus_input_offset_3_2;
  delay_66_q_net <= pixel_bus_input_offset_3_3;
  delay_68_q_net <= pixel_bus_input_offset_3_4;
  delay_70_q_net <= pixel_bus_input_offset_3_5;
  delay_50_q_net <= pixel_bus_input_offset_3_6;
  delay_52_q_net <= pixel_bus_input_offset_3_7;
  delay_54_q_net <= pixel_bus_input_offset_3_8;
  delay_63_q_net <= pixel_bus_input_offset_3_9;
  delay_56_q_net <= pixel_bus_input_offset_3_10;
  delay_58_q_net <= pixel_bus_input_offset_3_11;
  delay_61_q_net <= pixel_bus_input_offset_3_12;
  delay_84_q_net <= pixel_bus_input_offset_4_2;
  delay_90_q_net <= pixel_bus_input_offset_4_3;
  delay_92_q_net <= pixel_bus_input_offset_4_4;
  delay_94_q_net <= pixel_bus_input_offset_4_5;
  delay_74_q_net <= pixel_bus_input_offset_4_6;
  delay_76_q_net <= pixel_bus_input_offset_4_7;
  delay_78_q_net <= pixel_bus_input_offset_4_8;
  delay_87_q_net <= pixel_bus_input_offset_4_9;
  delay_80_q_net <= pixel_bus_input_offset_4_10;
  delay_82_q_net <= pixel_bus_input_offset_4_11;
  delay_85_q_net <= pixel_bus_input_offset_4_12;
  delay_3_q_net <= weight_bus_input_2;
  delay_5_q_net <= weight_bus_input_3;
  delay_7_q_net <= weight_bus_input_4;
  delay_9_q_net <= weight_bus_input_5;
  delay_11_q_net <= weight_bus_input_6;
  delay_13_q_net <= weight_bus_input_7;
  delay_15_q_net <= weight_bus_input_8;
  delay_24_q_net <= weight_bus_input_9;
  delay_17_q_net <= weight_bus_input_10;
  delay_19_q_net <= weight_bus_input_11;
  delay_21_q_net <= weight_bus_input_12;
  delay_25_q_net <= weight_bus_input_13;
  delay_41_q_net <= weight_bus_input_14;
  delay_43_q_net <= weight_bus_input_15;
  delay_45_q_net <= weight_bus_input_16;
  delay_47_q_net <= weight_bus_input_17;
  delay_27_q_net <= weight_bus_input_18;
  delay_29_q_net <= weight_bus_input_19;
  delay_31_q_net <= weight_bus_input_20;
  delay_40_q_net <= weight_bus_input_21;
  delay_33_q_net <= weight_bus_input_22;
  delay_35_q_net <= weight_bus_input_23;
  delay_38_q_net <= weight_bus_input_24;
  delay_49_q_net <= weight_bus_input_25;
  delay_65_q_net <= weight_bus_input_26;
  delay_67_q_net <= weight_bus_input_27;
  delay_69_q_net <= weight_bus_input_28;
  delay_71_q_net <= weight_bus_input_29;
  delay_51_q_net <= weight_bus_input_30;
  delay_53_q_net <= weight_bus_input_31;
  delay_55_q_net <= weight_bus_input_32;
  delay_64_q_net <= weight_bus_input_33;
  delay_57_q_net <= weight_bus_input_34;
  delay_59_q_net <= weight_bus_input_35;
  delay_62_q_net <= weight_bus_input_36;
  delay_73_q_net <= weight_bus_input_37;
  delay_89_q_net <= weight_bus_input_38;
  delay_91_q_net <= weight_bus_input_39;
  delay_93_q_net <= weight_bus_input_40;
  delay_95_q_net <= weight_bus_input_41;
  delay_75_q_net <= weight_bus_input_42;
  delay_77_q_net <= weight_bus_input_43;
  delay_79_q_net <= weight_bus_input_44;
  delay_88_q_net <= weight_bus_input_45;
  delay_81_q_net <= weight_bus_input_46;
  delay_83_q_net <= weight_bus_input_47;
  delay_86_q_net <= weight_bus_input_48;
  delay_97_q_net <= weight_bus_input_49;
  delay_113_q_net <= weight_bus_input_50;
  delay_115_q_net <= weight_bus_input_51;
  delay_117_q_net <= weight_bus_input_52;
  delay_119_q_net <= weight_bus_input_53;
  delay_99_q_net <= weight_bus_input_54;
  delay_101_q_net <= weight_bus_input_55;
  delay_103_q_net <= weight_bus_input_56;
  delay_112_q_net <= weight_bus_input_57;
  delay_105_q_net <= weight_bus_input_58;
  delay_107_q_net <= weight_bus_input_59;
  delay_110_q_net <= weight_bus_input_60;
  last_out_q_net <= weight_bus_input_61;
  enable_passthrough_case_0_y_net <= valid_bus_input_2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  accumlator_kernel_results : entity xil_defaultlib.mh_accumlator_kernel_results_x8 
  port map (
    slice_input_0 => accumulator_0_q_net_x3,
    slice_enable_0 => delay2_q_net_x3,
    slice_input_1 => accumulator_0_q_net_x2,
    slice_enable_1 => delay2_q_net_x2,
    slice_input_2 => accumulator_0_q_net_x1,
    slice_enable_2 => delay2_q_net_x1,
    slice_input_3 => accumulator_0_q_net_x0,
    slice_enable_3 => delay2_q_net_x0,
    slice_input_4 => accumulator_0_q_net,
    slice_enable_4 => delay2_q_net,
    reset_collector => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net
  );
  accumulator_offset_0 : entity xil_defaultlib.mh_accumulator_offset_0_x8 
  port map (
    input_value => last_combine_s_net_x3,
    input_valid => delay_addition4_q_net_x3,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x3,
    accumulator_valid => delay2_q_net_x3
  );
  accumulator_offset_1 : entity xil_defaultlib.mh_accumulator_offset_1_x8 
  port map (
    input_value => last_combine_s_net_x2,
    input_valid => delay_addition4_q_net_x2,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x2,
    accumulator_valid => delay2_q_net_x2
  );
  accumulator_offset_2 : entity xil_defaultlib.mh_accumulator_offset_2_x8 
  port map (
    input_value => last_combine_s_net_x1,
    input_valid => delay_addition4_q_net_x1,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x1,
    accumulator_valid => delay2_q_net_x1
  );
  accumulator_offset_3 : entity xil_defaultlib.mh_accumulator_offset_3_x8 
  port map (
    input_value => last_combine_s_net_x0,
    input_valid => delay_addition4_q_net_x0,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net_x0,
    accumulator_valid => delay2_q_net_x0
  );
  accumulator_offset_4 : entity xil_defaultlib.mh_accumulator_offset_4_x8 
  port map (
    input_value => last_combine_s_net,
    input_valid => delay_addition4_q_net,
    last_row => delay_addition4_q_net_x4,
    hard_reset => delay_addition8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    accumulator_output => accumulator_0_q_net,
    accumulator_valid => delay2_q_net
  );
  multiple_and_add_offset_0 : entity xil_defaultlib.mh_multiple_and_add_offset_0_x8 
  port map (
    pixel_0 => delay_96_q_net,
    weight_0 => delay_1_q_net,
    pixel_1 => delay_108_q_net,
    weight_1 => delay_3_q_net,
    pixel_2 => delay_114_q_net,
    weight_2 => delay_5_q_net,
    pixel_3 => delay_116_q_net,
    weight_3 => delay_7_q_net,
    pixel_4 => delay_118_q_net,
    weight_4 => delay_9_q_net,
    pixel_5 => delay_98_q_net,
    weight_5 => delay_11_q_net,
    pixel_6 => delay_100_q_net,
    weight_6 => delay_13_q_net,
    pixel_7 => delay_102_q_net,
    weight_7 => delay_15_q_net,
    pixel_8 => delay_111_q_net,
    weight_8 => delay_24_q_net,
    pixel_9 => delay_104_q_net,
    weight_9 => delay_17_q_net,
    pixel_10 => delay_106_q_net,
    weight_10 => delay_19_q_net,
    pixel_11 => delay_109_q_net,
    weight_11 => delay_21_q_net,
    valid_data => enable_passthrough_case_1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x3,
    valid_out => delay_addition4_q_net_x3
  );
  multiple_and_add_offset_1 : entity xil_defaultlib.mh_multiple_and_add_offset_1_x8 
  port map (
    pixel_0 => delay_0_q_net,
    weight_0 => delay_25_q_net,
    pixel_1 => delay_2_q_net,
    weight_1 => delay_41_q_net,
    pixel_2 => delay_4_q_net,
    weight_2 => delay_43_q_net,
    pixel_3 => delay_6_q_net,
    weight_3 => delay_45_q_net,
    pixel_4 => delay_8_q_net,
    weight_4 => delay_47_q_net,
    pixel_5 => delay_10_q_net,
    weight_5 => delay_27_q_net,
    pixel_6 => delay_12_q_net,
    weight_6 => delay_29_q_net,
    pixel_7 => delay_14_q_net,
    weight_7 => delay_31_q_net,
    pixel_8 => delay_23_q_net,
    weight_8 => delay_40_q_net,
    pixel_9 => delay_16_q_net,
    weight_9 => delay_33_q_net,
    pixel_10 => delay_18_q_net,
    weight_10 => delay_35_q_net,
    pixel_11 => delay_20_q_net,
    weight_11 => delay_38_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x2,
    valid_out => delay_addition4_q_net_x2
  );
  multiple_and_add_offset_2 : entity xil_defaultlib.mh_multiple_and_add_offset_2_x8 
  port map (
    pixel_0 => delay_22_q_net,
    weight_0 => delay_49_q_net,
    pixel_1 => delay_36_q_net,
    weight_1 => delay_65_q_net,
    pixel_2 => delay_42_q_net,
    weight_2 => delay_67_q_net,
    pixel_3 => delay_44_q_net,
    weight_3 => delay_69_q_net,
    pixel_4 => delay_46_q_net,
    weight_4 => delay_71_q_net,
    pixel_5 => delay_26_q_net,
    weight_5 => delay_51_q_net,
    pixel_6 => delay_28_q_net,
    weight_6 => delay_53_q_net,
    pixel_7 => delay_30_q_net,
    weight_7 => delay_55_q_net,
    pixel_8 => delay_39_q_net,
    weight_8 => delay_64_q_net,
    pixel_9 => delay_32_q_net,
    weight_9 => delay_57_q_net,
    pixel_10 => delay_34_q_net,
    weight_10 => delay_59_q_net,
    pixel_11 => delay_37_q_net,
    weight_11 => delay_62_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x1,
    valid_out => delay_addition4_q_net_x1
  );
  multiple_and_add_offset_3 : entity xil_defaultlib.mh_multiple_and_add_offset_3_x8 
  port map (
    pixel_0 => delay_48_q_net,
    weight_0 => delay_73_q_net,
    pixel_1 => delay_60_q_net,
    weight_1 => delay_89_q_net,
    pixel_2 => delay_66_q_net,
    weight_2 => delay_91_q_net,
    pixel_3 => delay_68_q_net,
    weight_3 => delay_93_q_net,
    pixel_4 => delay_70_q_net,
    weight_4 => delay_95_q_net,
    pixel_5 => delay_50_q_net,
    weight_5 => delay_75_q_net,
    pixel_6 => delay_52_q_net,
    weight_6 => delay_77_q_net,
    pixel_7 => delay_54_q_net,
    weight_7 => delay_79_q_net,
    pixel_8 => delay_63_q_net,
    weight_8 => delay_88_q_net,
    pixel_9 => delay_56_q_net,
    weight_9 => delay_81_q_net,
    pixel_10 => delay_58_q_net,
    weight_10 => delay_83_q_net,
    pixel_11 => delay_61_q_net,
    weight_11 => delay_86_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net_x0,
    valid_out => delay_addition4_q_net_x0
  );
  multiple_and_add_offset_4 : entity xil_defaultlib.mh_multiple_and_add_offset_4_x8 
  port map (
    pixel_0 => delay_72_q_net,
    weight_0 => delay_97_q_net,
    pixel_1 => delay_84_q_net,
    weight_1 => delay_113_q_net,
    pixel_2 => delay_90_q_net,
    weight_2 => delay_115_q_net,
    pixel_3 => delay_92_q_net,
    weight_3 => delay_117_q_net,
    pixel_4 => delay_94_q_net,
    weight_4 => delay_119_q_net,
    pixel_5 => delay_74_q_net,
    weight_5 => delay_99_q_net,
    pixel_6 => delay_76_q_net,
    weight_6 => delay_101_q_net,
    pixel_7 => delay_78_q_net,
    weight_7 => delay_103_q_net,
    pixel_8 => delay_87_q_net,
    weight_8 => delay_112_q_net,
    pixel_9 => delay_80_q_net,
    weight_9 => delay_105_q_net,
    pixel_10 => delay_82_q_net,
    weight_10 => delay_107_q_net,
    pixel_11 => delay_85_q_net,
    weight_11 => delay_110_q_net,
    valid_data => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    slice_out => last_combine_s_net,
    valid_out => delay_addition4_q_net
  );
  delay_addition_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_1_q_net
  );
  delay_addition_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition_2_q_net
  );
  delay_addition1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => last_out_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition1_q_net
  );
  delay_addition2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition2_q_net
  );
  delay_addition3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition3_q_net
  );
  delay_addition4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition4_q_net_x4
  );
  delay_addition5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition5_q_net
  );
  delay_addition6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition6_q_net
  );
  delay_addition7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition7_q_net
  );
  delay_addition8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_addition7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_addition8_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math/Subsystem
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_subsystem is
  port (
    kernel_result_0 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_0 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_1 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_1 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_2 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_2 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_3 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_3 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_4 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_4 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_5 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_5 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_6 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_6 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_7 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_7 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_8 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_8 : in std_logic_vector( 1-1 downto 0 );
    kernel_result_9 : in std_logic_vector( 128-1 downto 0 );
    kernel_result_valid_9 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_result_output : out std_logic_vector( 128-1 downto 0 );
    kernel_result_output_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_result_array_position : out std_logic_vector( 12-1 downto 0 );
    kernel_result_row_depth_position : out std_logic_vector( 12-1 downto 0 );
    finished_cube : out std_logic_vector( 1-1 downto 0 )
  );
end mh_subsystem;
architecture structural of mh_subsystem is 
  signal mux_enable_delay_8_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_enable_delay_9_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_enable_delay_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_enable_delay_5_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_1_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_enable_delay_7_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_0_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_enable_delay_6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_slice_4_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_8_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_9_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_5_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_7_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_2_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_6_y_net : std_logic_vector( 128-1 downto 0 );
  signal mux_slice_3_y_net : std_logic_vector( 128-1 downto 0 );
  signal output_or_block_y_net : std_logic_vector( 128-1 downto 0 );
  signal kernel_result_array_offset_op_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x0 : std_logic_vector( 128-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x7 : std_logic_vector( 128-1 downto 0 );
  signal kernel_result_array_offset1_op_net : std_logic_vector( 12-1 downto 0 );
  signal delay_enable_4_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x5 : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal accumulator_kernel_result_0_q_net_x1 : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x6 : std_logic_vector( 128-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x4 : std_logic_vector( 128-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x2 : std_logic_vector( 128-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_enable_4_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal output_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal base_value_op_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x8 : std_logic_vector( 128-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x3 : std_logic_vector( 128-1 downto 0 );
  signal max_value_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_enable_delay_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_enable_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_enable_delay_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 12-1 downto 0 );
  signal mux_enable_delay_3_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 32-1 downto 0 );
begin
  kernel_result_output <= output_or_block_y_net;
  kernel_result_output_valid <= output_enable_y_net;
  kernel_result_array_position <= kernel_result_array_offset_op_net;
  kernel_result_row_depth_position <= kernel_result_array_offset1_op_net;
  finished_cube <= switch_to_zero_y_net;
  accumulator_kernel_result_0_q_net_x8 <= kernel_result_0;
  delay_enable_4_q_net_x8 <= kernel_result_valid_0;
  accumulator_kernel_result_0_q_net_x7 <= kernel_result_1;
  delay_enable_4_q_net_x7 <= kernel_result_valid_1;
  accumulator_kernel_result_0_q_net_x6 <= kernel_result_2;
  delay_enable_4_q_net_x6 <= kernel_result_valid_2;
  accumulator_kernel_result_0_q_net_x5 <= kernel_result_3;
  delay_enable_4_q_net_x5 <= kernel_result_valid_3;
  accumulator_kernel_result_0_q_net_x4 <= kernel_result_4;
  delay_enable_4_q_net_x4 <= kernel_result_valid_4;
  accumulator_kernel_result_0_q_net_x3 <= kernel_result_5;
  delay_enable_4_q_net_x3 <= kernel_result_valid_5;
  accumulator_kernel_result_0_q_net_x2 <= kernel_result_6;
  delay_enable_4_q_net_x2 <= kernel_result_valid_6;
  accumulator_kernel_result_0_q_net_x1 <= kernel_result_7;
  delay_enable_4_q_net_x1 <= kernel_result_valid_7;
  accumulator_kernel_result_0_q_net_x0 <= kernel_result_8;
  delay_enable_4_q_net_x0 <= kernel_result_valid_8;
  accumulator_kernel_result_0_q_net <= kernel_result_9;
  delay_enable_4_q_net <= kernel_result_valid_9;
  clk_net <= clk_1;
  ce_net <= ce_1;
  base_value : entity xil_defaultlib.sysgen_relational_7b3bb090a4 
  port map (
    clr => '0',
    a => kernel_result_array_offset_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => base_value_op_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_70e8a7b61d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_162ea2571e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => max_value_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  kernel_result_array_offset : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 1095,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i3",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 12
  )
  port map (
    rst => "0",
    clr => '0',
    en => output_enable_y_net,
    clk => clk_net,
    ce => ce_net,
    op => kernel_result_array_offset_op_net
  );
  kernel_result_array_offset1 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 1095,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i3",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 12
  )
  port map (
    rst => "0",
    clr => '0',
    en => switch_to_zero_y_net,
    clk => clk_net,
    ce => ce_net,
    op => kernel_result_array_offset1_op_net
  );
  mux_enable_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_0_q_net
  );
  mux_enable_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_1_q_net
  );
  mux_enable_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_2_q_net
  );
  mux_enable_delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_3_q_net
  );
  mux_enable_delay_4 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_4_q_net
  );
  mux_enable_delay_5 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_5_q_net
  );
  mux_enable_delay_6 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_6_q_net
  );
  mux_enable_delay_7 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_7_q_net
  );
  mux_enable_delay_8 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_8_q_net
  );
  mux_enable_delay_9 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_enable_4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_9_q_net
  );
  max_value : entity xil_defaultlib.sysgen_relational_75c30532cf 
  port map (
    clr => '0',
    a => kernel_result_array_offset_op_net,
    b => constant3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => max_value_op_net
  );
  mux_slice_0 : entity xil_defaultlib.sysgen_mux_57d8a3c9d4 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x8,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x8,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_0_y_net
  );
  mux_slice_1 : entity xil_defaultlib.sysgen_mux_d116dd3dfc 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x7,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x7,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_1_y_net
  );
  mux_slice_2 : entity xil_defaultlib.sysgen_mux_67eb8c2e6f 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x6,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x6,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_2_y_net
  );
  mux_slice_3 : entity xil_defaultlib.sysgen_mux_5fa8cfdba3 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x5,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_3_y_net
  );
  mux_slice_4 : entity xil_defaultlib.sysgen_mux_53b009d61b 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x4,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_4_y_net
  );
  mux_slice_5 : entity xil_defaultlib.sysgen_mux_57d8a3c9d4 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x3,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_5_y_net
  );
  mux_slice_6 : entity xil_defaultlib.sysgen_mux_d116dd3dfc 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x2,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_6_y_net
  );
  mux_slice_7 : entity xil_defaultlib.sysgen_mux_67eb8c2e6f 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x1,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_7_y_net
  );
  mux_slice_8 : entity xil_defaultlib.sysgen_mux_5fa8cfdba3 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net_x0,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_8_y_net
  );
  mux_slice_9 : entity xil_defaultlib.sysgen_mux_53b009d61b 
  port map (
    clr => '0',
    sel => delay_enable_4_q_net,
    d0 => constant1_op_net,
    d1 => accumulator_kernel_result_0_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_slice_9_y_net
  );
  output_enable : entity xil_defaultlib.sysgen_logical_c7239c6e66 
  port map (
    clr => '0',
    d0 => mux_enable_delay_0_q_net,
    d1 => mux_enable_delay_1_q_net,
    d2 => mux_enable_delay_2_q_net,
    d3 => mux_enable_delay_3_q_net,
    d4 => mux_enable_delay_4_q_net,
    d5 => mux_enable_delay_5_q_net,
    d6 => mux_enable_delay_6_q_net,
    d7 => mux_enable_delay_7_q_net,
    d8 => mux_enable_delay_8_q_net,
    d9 => mux_enable_delay_9_q_net,
    clk => clk_net,
    ce => ce_net,
    y => output_enable_y_net
  );
  output_or_block : entity xil_defaultlib.sysgen_logical_b33b7318c8 
  port map (
    clr => '0',
    d0 => mux_slice_0_y_net,
    d1 => mux_slice_1_y_net,
    d2 => mux_slice_2_y_net,
    d3 => mux_slice_3_y_net,
    d4 => mux_slice_4_y_net,
    d5 => mux_slice_5_y_net,
    d6 => mux_slice_6_y_net,
    d7 => mux_slice_7_y_net,
    d8 => mux_slice_8_y_net,
    d9 => mux_slice_9_y_net,
    clk => clk_net,
    ce => ce_net,
    y => output_or_block_y_net
  );
  switch_to_zero : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => base_value_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => switch_to_zero_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Math
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_math is
  port (
    in_pixel_0_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_0 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_1 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_2 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_3 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_0_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_1_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_2_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_3_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_4_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_5_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_6_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_7_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_8_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_9_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_10_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_pixel_11_at_offset_4 : in std_logic_vector( 12-1 downto 0 );
    in_weight_0_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_0 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_1 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_2 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_3 : in std_logic_vector( 18-1 downto 0 );
    in_weight_0_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_1_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_2_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_3_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_4_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_5_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_6_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_7_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_8_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_9_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_10_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    in_weight_11_at_offset_4 : in std_logic_vector( 18-1 downto 0 );
    valid_data_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_output : out std_logic_vector( 128-1 downto 0 );
    valid_kernel_output : out std_logic_vector( 1-1 downto 0 );
    kernel_result_array_position : out std_logic_vector( 12-1 downto 0 );
    kernel_result_row_depth_position : out std_logic_vector( 12-1 downto 0 )
  );
end mh_math;
architecture structural of mh_math is 
  signal x12_bit_bin_value_0_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal output_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal kernel_result_array_offset1_op_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal kernel_result_array_offset_op_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal output_or_block_y_net : std_logic_vector( 128-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x3 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_0_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_22_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal delay_14_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_36_q_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_96_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_4_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_10_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_12_q_net : std_logic_vector( 12-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_16_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_18_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_72_q_net : std_logic_vector( 12-1 downto 0 );
  signal data_valid_out_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal delay_20_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_42_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_23_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_44_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_46_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_6_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_26_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_28_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_30_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_48_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_39_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_47_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_27_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_40_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_33_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_31_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_61_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_74_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_111_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_49_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_38_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_68_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_24_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_32_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_65_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_82_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_67_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_98_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_29_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_108_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_69_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_80_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_54_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_85_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_114_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_52_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_37_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_17_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_100_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_45_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_71_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_50_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_78_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_60_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_94_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_56_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_76_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_70_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_63_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_87_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_116_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_84_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_102_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_106_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_109_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_104_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_34_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_92_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_58_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_118_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_90_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_25_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_66_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay_41_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_43_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x0 : std_logic_vector( 128-1 downto 0 );
  signal enable_passthrough_case_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x1 : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x5 : std_logic_vector( 128-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal delay_81_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_53_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_57_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_83_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_115_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_64_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_95_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_117_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_112_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal delay_79_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_75_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_86_q_net : std_logic_vector( 18-1 downto 0 );
  signal switch_to_zero_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_55_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_enable_4_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x2 : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_99_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_110_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x3 : std_logic_vector( 128-1 downto 0 );
  signal delay_105_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_59_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_kernel_result_0_q_net : std_logic_vector( 128-1 downto 0 );
  signal delay_enable_4_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x7 : std_logic_vector( 128-1 downto 0 );
  signal delay_101_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_1_y_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_91_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_enable_4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal last_out_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_93_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_51_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_113_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x8 : std_logic_vector( 128-1 downto 0 );
  signal delay_119_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_97_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_62_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_89_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_107_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_73_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_88_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x6 : std_logic_vector( 128-1 downto 0 );
  signal delay_77_q_net : std_logic_vector( 18-1 downto 0 );
  signal accumulator_kernel_result_0_q_net_x4 : std_logic_vector( 128-1 downto 0 );
  signal delay_103_q_net : std_logic_vector( 18-1 downto 0 );
  signal enable_passthrough_case_0_y_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay_enable_4_q_net_x3 : std_logic_vector( 1-1 downto 0 );
begin
  kernel_output <= output_or_block_y_net;
  valid_kernel_output <= output_enable_y_net;
  kernel_result_array_position <= kernel_result_array_offset_op_net;
  kernel_result_row_depth_position <= kernel_result_array_offset1_op_net;
  x12_bit_bin_value_0_q_net_x8 <= in_pixel_0_at_offset_0;
  x12_bit_bin_value_1_q_net_x8 <= in_pixel_1_at_offset_0;
  x12_bit_bin_value_2_q_net_x7 <= in_pixel_2_at_offset_0;
  x12_bit_bin_value_3_q_net_x8 <= in_pixel_3_at_offset_0;
  x12_bit_bin_value_4_q_net_x8 <= in_pixel_4_at_offset_0;
  x12_bit_bin_value_5_q_net_x8 <= in_pixel_5_at_offset_0;
  x12_bit_bin_value_6_q_net_x8 <= in_pixel_6_at_offset_0;
  x12_bit_bin_value_7_q_net_x8 <= in_pixel_7_at_offset_0;
  x12_bit_bin_value_8_q_net_x8 <= in_pixel_8_at_offset_0;
  x12_bit_bin_value_9_q_net_x8 <= in_pixel_9_at_offset_0;
  x12_bit_bin_value_10_q_net_x8 <= in_pixel_10_at_offset_0;
  x12_bit_bin_value_11_q_net_x8 <= in_pixel_11_at_offset_0;
  x12_bit_bin_value_0_q_net_x7 <= in_pixel_0_at_offset_1;
  x12_bit_bin_value_1_q_net_x7 <= in_pixel_1_at_offset_1;
  x12_bit_bin_value_2_q_net_x6 <= in_pixel_2_at_offset_1;
  x12_bit_bin_value_3_q_net_x7 <= in_pixel_3_at_offset_1;
  x12_bit_bin_value_4_q_net_x7 <= in_pixel_4_at_offset_1;
  x12_bit_bin_value_5_q_net_x7 <= in_pixel_5_at_offset_1;
  x12_bit_bin_value_6_q_net_x7 <= in_pixel_6_at_offset_1;
  x12_bit_bin_value_7_q_net_x7 <= in_pixel_7_at_offset_1;
  x12_bit_bin_value_8_q_net_x7 <= in_pixel_8_at_offset_1;
  x12_bit_bin_value_9_q_net_x7 <= in_pixel_9_at_offset_1;
  x12_bit_bin_value_10_q_net_x7 <= in_pixel_10_at_offset_1;
  x12_bit_bin_value_11_q_net_x7 <= in_pixel_11_at_offset_1;
  x12_bit_bin_value_0_q_net_x6 <= in_pixel_0_at_offset_2;
  x12_bit_bin_value_1_q_net_x6 <= in_pixel_1_at_offset_2;
  x12_bit_bin_value_2_q_net_x5 <= in_pixel_2_at_offset_2;
  x12_bit_bin_value_3_q_net_x6 <= in_pixel_3_at_offset_2;
  x12_bit_bin_value_4_q_net_x6 <= in_pixel_4_at_offset_2;
  x12_bit_bin_value_5_q_net_x6 <= in_pixel_5_at_offset_2;
  x12_bit_bin_value_6_q_net_x6 <= in_pixel_6_at_offset_2;
  x12_bit_bin_value_7_q_net_x6 <= in_pixel_7_at_offset_2;
  x12_bit_bin_value_8_q_net_x6 <= in_pixel_8_at_offset_2;
  x12_bit_bin_value_9_q_net_x6 <= in_pixel_9_at_offset_2;
  x12_bit_bin_value_10_q_net_x6 <= in_pixel_10_at_offset_2;
  x12_bit_bin_value_11_q_net_x6 <= in_pixel_11_at_offset_2;
  x12_bit_bin_value_0_q_net_x5 <= in_pixel_0_at_offset_3;
  x12_bit_bin_value_1_q_net_x5 <= in_pixel_1_at_offset_3;
  x12_bit_bin_value_2_q_net_x8 <= in_pixel_2_at_offset_3;
  x12_bit_bin_value_3_q_net_x5 <= in_pixel_3_at_offset_3;
  x12_bit_bin_value_4_q_net_x5 <= in_pixel_4_at_offset_3;
  x12_bit_bin_value_5_q_net_x5 <= in_pixel_5_at_offset_3;
  x12_bit_bin_value_6_q_net_x5 <= in_pixel_6_at_offset_3;
  x12_bit_bin_value_7_q_net_x4 <= in_pixel_7_at_offset_3;
  x12_bit_bin_value_8_q_net_x5 <= in_pixel_8_at_offset_3;
  x12_bit_bin_value_9_q_net_x5 <= in_pixel_9_at_offset_3;
  x12_bit_bin_value_10_q_net_x5 <= in_pixel_10_at_offset_3;
  x12_bit_bin_value_11_q_net_x5 <= in_pixel_11_at_offset_3;
  x12_bit_bin_value_0_q_net_x4 <= in_pixel_0_at_offset_4;
  x12_bit_bin_value_1_q_net_x4 <= in_pixel_1_at_offset_4;
  x12_bit_bin_value_2_q_net_x4 <= in_pixel_2_at_offset_4;
  x12_bit_bin_value_3_q_net_x4 <= in_pixel_3_at_offset_4;
  x12_bit_bin_value_4_q_net_x4 <= in_pixel_4_at_offset_4;
  x12_bit_bin_value_5_q_net_x4 <= in_pixel_5_at_offset_4;
  x12_bit_bin_value_6_q_net_x4 <= in_pixel_6_at_offset_4;
  x12_bit_bin_value_7_q_net_x3 <= in_pixel_7_at_offset_4;
  x12_bit_bin_value_8_q_net_x4 <= in_pixel_8_at_offset_4;
  x12_bit_bin_value_9_q_net_x4 <= in_pixel_9_at_offset_4;
  x12_bit_bin_value_10_q_net_x4 <= in_pixel_10_at_offset_4;
  x12_bit_bin_value_11_q_net_x4 <= in_pixel_11_at_offset_4;
  x12_bit_bin_value_0_q_net_x3 <= in_weight_0_at_offset_0;
  x12_bit_bin_value_1_q_net_x3 <= in_weight_1_at_offset_0;
  x12_bit_bin_value_2_q_net_x3 <= in_weight_2_at_offset_0;
  x12_bit_bin_value_3_q_net_x3 <= in_weight_3_at_offset_0;
  x12_bit_bin_value_4_q_net_x3 <= in_weight_4_at_offset_0;
  x12_bit_bin_value_5_q_net_x3 <= in_weight_5_at_offset_0;
  x12_bit_bin_value_6_q_net_x3 <= in_weight_6_at_offset_0;
  x12_bit_bin_value_7_q_net_x2 <= in_weight_7_at_offset_0;
  x12_bit_bin_value_8_q_net_x3 <= in_weight_8_at_offset_0;
  x12_bit_bin_value_9_q_net_x3 <= in_weight_9_at_offset_0;
  x12_bit_bin_value_10_q_net_x3 <= in_weight_10_at_offset_0;
  x12_bit_bin_value_11_q_net_x3 <= in_weight_11_at_offset_0;
  x12_bit_bin_value_0_q_net_x2 <= in_weight_0_at_offset_1;
  x12_bit_bin_value_1_q_net_x2 <= in_weight_1_at_offset_1;
  x12_bit_bin_value_2_q_net_x2 <= in_weight_2_at_offset_1;
  x12_bit_bin_value_3_q_net_x2 <= in_weight_3_at_offset_1;
  x12_bit_bin_value_4_q_net_x2 <= in_weight_4_at_offset_1;
  x12_bit_bin_value_5_q_net_x2 <= in_weight_5_at_offset_1;
  x12_bit_bin_value_6_q_net_x2 <= in_weight_6_at_offset_1;
  x12_bit_bin_value_7_q_net_x1 <= in_weight_7_at_offset_1;
  x12_bit_bin_value_8_q_net_x2 <= in_weight_8_at_offset_1;
  x12_bit_bin_value_9_q_net_x2 <= in_weight_9_at_offset_1;
  x12_bit_bin_value_10_q_net_x2 <= in_weight_10_at_offset_1;
  x12_bit_bin_value_11_q_net_x2 <= in_weight_11_at_offset_1;
  x12_bit_bin_value_0_q_net_x1 <= in_weight_0_at_offset_2;
  x12_bit_bin_value_1_q_net_x1 <= in_weight_1_at_offset_2;
  x12_bit_bin_value_2_q_net_x1 <= in_weight_2_at_offset_2;
  x12_bit_bin_value_3_q_net_x1 <= in_weight_3_at_offset_2;
  x12_bit_bin_value_4_q_net_x1 <= in_weight_4_at_offset_2;
  x12_bit_bin_value_5_q_net_x1 <= in_weight_5_at_offset_2;
  x12_bit_bin_value_6_q_net_x1 <= in_weight_6_at_offset_2;
  x12_bit_bin_value_7_q_net_x5 <= in_weight_7_at_offset_2;
  x12_bit_bin_value_8_q_net_x1 <= in_weight_8_at_offset_2;
  x12_bit_bin_value_9_q_net_x1 <= in_weight_9_at_offset_2;
  x12_bit_bin_value_10_q_net_x1 <= in_weight_10_at_offset_2;
  x12_bit_bin_value_11_q_net_x1 <= in_weight_11_at_offset_2;
  x12_bit_bin_value_0_q_net_x0 <= in_weight_0_at_offset_3;
  x12_bit_bin_value_1_q_net_x0 <= in_weight_1_at_offset_3;
  x12_bit_bin_value_2_q_net_x0 <= in_weight_2_at_offset_3;
  x12_bit_bin_value_3_q_net_x0 <= in_weight_3_at_offset_3;
  x12_bit_bin_value_4_q_net_x0 <= in_weight_4_at_offset_3;
  x12_bit_bin_value_5_q_net_x0 <= in_weight_5_at_offset_3;
  x12_bit_bin_value_6_q_net_x0 <= in_weight_6_at_offset_3;
  x12_bit_bin_value_7_q_net_x0 <= in_weight_7_at_offset_3;
  x12_bit_bin_value_8_q_net_x0 <= in_weight_8_at_offset_3;
  x12_bit_bin_value_9_q_net_x0 <= in_weight_9_at_offset_3;
  x12_bit_bin_value_10_q_net_x0 <= in_weight_10_at_offset_3;
  x12_bit_bin_value_11_q_net_x0 <= in_weight_11_at_offset_3;
  x12_bit_bin_value_0_q_net <= in_weight_0_at_offset_4;
  x12_bit_bin_value_1_q_net <= in_weight_1_at_offset_4;
  x12_bit_bin_value_2_q_net <= in_weight_2_at_offset_4;
  x12_bit_bin_value_3_q_net <= in_weight_3_at_offset_4;
  x12_bit_bin_value_4_q_net <= in_weight_4_at_offset_4;
  x12_bit_bin_value_5_q_net <= in_weight_5_at_offset_4;
  x12_bit_bin_value_6_q_net <= in_weight_6_at_offset_4;
  x12_bit_bin_value_7_q_net <= in_weight_7_at_offset_4;
  x12_bit_bin_value_8_q_net <= in_weight_8_at_offset_4;
  x12_bit_bin_value_9_q_net <= in_weight_9_at_offset_4;
  x12_bit_bin_value_10_q_net <= in_weight_10_at_offset_4;
  x12_bit_bin_value_11_q_net <= in_weight_11_at_offset_4;
  data_valid_out_delay_q_net <= valid_data_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  kernel_organizer : entity xil_defaultlib.mh_kernel_organizer 
  port map (
    in_pixel_0_at_offset_0 => x12_bit_bin_value_0_q_net_x8,
    in_pixel_1_at_offset_0 => x12_bit_bin_value_1_q_net_x8,
    in_pixel_2_at_offset_0 => x12_bit_bin_value_2_q_net_x7,
    in_pixel_3_at_offset_0 => x12_bit_bin_value_3_q_net_x8,
    in_pixel_4_at_offset_0 => x12_bit_bin_value_4_q_net_x8,
    in_pixel_5_at_offset_0 => x12_bit_bin_value_5_q_net_x8,
    in_pixel_6_at_offset_0 => x12_bit_bin_value_6_q_net_x8,
    in_pixel_7_at_offset_0 => x12_bit_bin_value_7_q_net_x8,
    in_pixel_8_at_offset_0 => x12_bit_bin_value_8_q_net_x8,
    in_pixel_9_at_offset_0 => x12_bit_bin_value_9_q_net_x8,
    in_pixel_10_at_offset_0 => x12_bit_bin_value_10_q_net_x8,
    in_pixel_11_at_offset_0 => x12_bit_bin_value_11_q_net_x8,
    in_pixel_0_at_offset_1 => x12_bit_bin_value_0_q_net_x7,
    in_pixel_1_at_offset_1 => x12_bit_bin_value_1_q_net_x7,
    in_pixel_2_at_offset_1 => x12_bit_bin_value_2_q_net_x6,
    in_pixel_3_at_offset_1 => x12_bit_bin_value_3_q_net_x7,
    in_pixel_4_at_offset_1 => x12_bit_bin_value_4_q_net_x7,
    in_pixel_5_at_offset_1 => x12_bit_bin_value_5_q_net_x7,
    in_pixel_6_at_offset_1 => x12_bit_bin_value_6_q_net_x7,
    in_pixel_7_at_offset_1 => x12_bit_bin_value_7_q_net_x7,
    in_pixel_8_at_offset_1 => x12_bit_bin_value_8_q_net_x7,
    in_pixel_9_at_offset_1 => x12_bit_bin_value_9_q_net_x7,
    in_pixel_10_at_offset_1 => x12_bit_bin_value_10_q_net_x7,
    in_pixel_11_at_offset_1 => x12_bit_bin_value_11_q_net_x7,
    in_pixel_0_at_offset_2 => x12_bit_bin_value_0_q_net_x6,
    in_pixel_1_at_offset_2 => x12_bit_bin_value_1_q_net_x6,
    in_pixel_2_at_offset_2 => x12_bit_bin_value_2_q_net_x5,
    in_pixel_3_at_offset_2 => x12_bit_bin_value_3_q_net_x6,
    in_pixel_4_at_offset_2 => x12_bit_bin_value_4_q_net_x6,
    in_pixel_5_at_offset_2 => x12_bit_bin_value_5_q_net_x6,
    in_pixel_6_at_offset_2 => x12_bit_bin_value_6_q_net_x6,
    in_pixel_7_at_offset_2 => x12_bit_bin_value_7_q_net_x6,
    in_pixel_8_at_offset_2 => x12_bit_bin_value_8_q_net_x6,
    in_pixel_9_at_offset_2 => x12_bit_bin_value_9_q_net_x6,
    in_pixel_10_at_offset_2 => x12_bit_bin_value_10_q_net_x6,
    in_pixel_11_at_offset_2 => x12_bit_bin_value_11_q_net_x6,
    in_pixel_0_at_offset_3 => x12_bit_bin_value_0_q_net_x5,
    in_pixel_1_at_offset_3 => x12_bit_bin_value_1_q_net_x5,
    in_pixel_2_at_offset_3 => x12_bit_bin_value_2_q_net_x8,
    in_pixel_3_at_offset_3 => x12_bit_bin_value_3_q_net_x5,
    in_pixel_4_at_offset_3 => x12_bit_bin_value_4_q_net_x5,
    in_pixel_5_at_offset_3 => x12_bit_bin_value_5_q_net_x5,
    in_pixel_6_at_offset_3 => x12_bit_bin_value_6_q_net_x5,
    in_pixel_7_at_offset_3 => x12_bit_bin_value_7_q_net_x4,
    in_pixel_8_at_offset_3 => x12_bit_bin_value_8_q_net_x5,
    in_pixel_9_at_offset_3 => x12_bit_bin_value_9_q_net_x5,
    in_pixel_10_at_offset_3 => x12_bit_bin_value_10_q_net_x5,
    in_pixel_11_at_offset_3 => x12_bit_bin_value_11_q_net_x5,
    in_pixel_0_at_offset_4 => x12_bit_bin_value_0_q_net_x4,
    in_pixel_1_at_offset_4 => x12_bit_bin_value_1_q_net_x4,
    in_pixel_2_at_offset_4 => x12_bit_bin_value_2_q_net_x4,
    in_pixel_3_at_offset_4 => x12_bit_bin_value_3_q_net_x4,
    in_pixel_4_at_offset_4 => x12_bit_bin_value_4_q_net_x4,
    in_pixel_5_at_offset_4 => x12_bit_bin_value_5_q_net_x4,
    in_pixel_6_at_offset_4 => x12_bit_bin_value_6_q_net_x4,
    in_pixel_7_at_offset_4 => x12_bit_bin_value_7_q_net_x3,
    in_pixel_8_at_offset_4 => x12_bit_bin_value_8_q_net_x4,
    in_pixel_9_at_offset_4 => x12_bit_bin_value_9_q_net_x4,
    in_pixel_10_at_offset_4 => x12_bit_bin_value_10_q_net_x4,
    in_pixel_11_at_offset_4 => x12_bit_bin_value_11_q_net_x4,
    in_weight_0_at_offset_0 => x12_bit_bin_value_0_q_net_x3,
    in_weight_1_at_offset_0 => x12_bit_bin_value_1_q_net_x3,
    in_weight_2_at_offset_0 => x12_bit_bin_value_2_q_net_x3,
    in_weight_3_at_offset_0 => x12_bit_bin_value_3_q_net_x3,
    in_weight_4_at_offset_0 => x12_bit_bin_value_4_q_net_x3,
    in_weight_5_at_offset_0 => x12_bit_bin_value_5_q_net_x3,
    in_weight_6_at_offset_0 => x12_bit_bin_value_6_q_net_x3,
    in_weight_7_at_offset_0 => x12_bit_bin_value_7_q_net_x2,
    in_weight_8_at_offset_0 => x12_bit_bin_value_8_q_net_x3,
    in_weight_9_at_offset_0 => x12_bit_bin_value_9_q_net_x3,
    in_weight_10_at_offset_0 => x12_bit_bin_value_10_q_net_x3,
    in_weight_11_at_offset_0 => x12_bit_bin_value_11_q_net_x3,
    in_weight_0_at_offset_1 => x12_bit_bin_value_0_q_net_x2,
    in_weight_1_at_offset_1 => x12_bit_bin_value_1_q_net_x2,
    in_weight_2_at_offset_1 => x12_bit_bin_value_2_q_net_x2,
    in_weight_3_at_offset_1 => x12_bit_bin_value_3_q_net_x2,
    in_weight_4_at_offset_1 => x12_bit_bin_value_4_q_net_x2,
    in_weight_5_at_offset_1 => x12_bit_bin_value_5_q_net_x2,
    in_weight_6_at_offset_1 => x12_bit_bin_value_6_q_net_x2,
    in_weight_7_at_offset_1 => x12_bit_bin_value_7_q_net_x1,
    in_weight_8_at_offset_1 => x12_bit_bin_value_8_q_net_x2,
    in_weight_9_at_offset_1 => x12_bit_bin_value_9_q_net_x2,
    in_weight_10_at_offset_1 => x12_bit_bin_value_10_q_net_x2,
    in_weight_11_at_offset_1 => x12_bit_bin_value_11_q_net_x2,
    in_weight_0_at_offset_2 => x12_bit_bin_value_0_q_net_x1,
    in_weight_1_at_offset_2 => x12_bit_bin_value_1_q_net_x1,
    in_weight_2_at_offset_2 => x12_bit_bin_value_2_q_net_x1,
    in_weight_3_at_offset_2 => x12_bit_bin_value_3_q_net_x1,
    in_weight_4_at_offset_2 => x12_bit_bin_value_4_q_net_x1,
    in_weight_5_at_offset_2 => x12_bit_bin_value_5_q_net_x1,
    in_weight_6_at_offset_2 => x12_bit_bin_value_6_q_net_x1,
    in_weight_7_at_offset_2 => x12_bit_bin_value_7_q_net_x5,
    in_weight_8_at_offset_2 => x12_bit_bin_value_8_q_net_x1,
    in_weight_9_at_offset_2 => x12_bit_bin_value_9_q_net_x1,
    in_weight_10_at_offset_2 => x12_bit_bin_value_10_q_net_x1,
    in_weight_11_at_offset_2 => x12_bit_bin_value_11_q_net_x1,
    in_weight_0_at_offset_3 => x12_bit_bin_value_0_q_net_x0,
    in_weight_1_at_offset_3 => x12_bit_bin_value_1_q_net_x0,
    in_weight_2_at_offset_3 => x12_bit_bin_value_2_q_net_x0,
    in_weight_3_at_offset_3 => x12_bit_bin_value_3_q_net_x0,
    in_weight_4_at_offset_3 => x12_bit_bin_value_4_q_net_x0,
    in_weight_5_at_offset_3 => x12_bit_bin_value_5_q_net_x0,
    in_weight_6_at_offset_3 => x12_bit_bin_value_6_q_net_x0,
    in_weight_7_at_offset_3 => x12_bit_bin_value_7_q_net_x0,
    in_weight_8_at_offset_3 => x12_bit_bin_value_8_q_net_x0,
    in_weight_9_at_offset_3 => x12_bit_bin_value_9_q_net_x0,
    in_weight_10_at_offset_3 => x12_bit_bin_value_10_q_net_x0,
    in_weight_11_at_offset_3 => x12_bit_bin_value_11_q_net_x0,
    in_weight_0_at_offset_4 => x12_bit_bin_value_0_q_net,
    in_weight_1_at_offset_4 => x12_bit_bin_value_1_q_net,
    in_weight_2_at_offset_4 => x12_bit_bin_value_2_q_net,
    in_weight_3_at_offset_4 => x12_bit_bin_value_3_q_net,
    in_weight_4_at_offset_4 => x12_bit_bin_value_4_q_net,
    in_weight_5_at_offset_4 => x12_bit_bin_value_5_q_net,
    in_weight_6_at_offset_4 => x12_bit_bin_value_6_q_net,
    in_weight_7_at_offset_4 => x12_bit_bin_value_7_q_net,
    in_weight_8_at_offset_4 => x12_bit_bin_value_8_q_net,
    in_weight_9_at_offset_4 => x12_bit_bin_value_9_q_net,
    in_weight_10_at_offset_4 => x12_bit_bin_value_10_q_net,
    in_weight_11_at_offset_4 => x12_bit_bin_value_11_q_net,
    valid_data_in => data_valid_out_delay_q_net,
    reset_to_known_state => switch_to_zero_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    pixel_group_offset_0_1 => delay_0_q_net,
    pixel_group_offset_1_1 => delay_22_q_net,
    pixel_group_offset_2_1 => delay_48_q_net,
    pixel_group_offset_3_1 => delay_72_q_net,
    pixel_group_offset_4_1 => delay_96_q_net,
    weights_1 => delay_1_q_net,
    kernel_result_valid_bus_0_1 => enable_passthrough_case_0_y_net_x7,
    kernel_result_valid_bus_1_1 => enable_passthrough_case_0_y_net_x6,
    kernel_result_valid_bus_2_1 => enable_passthrough_case_0_y_net_x5,
    kernel_result_valid_bus_3_1 => enable_passthrough_case_0_y_net_x4,
    kernel_result_valid_bus_4_1 => enable_passthrough_case_0_y_net_x3,
    kernel_result_valid_bus_5_1 => enable_passthrough_case_1_y_net_x3,
    kernel_result_valid_bus_6_1 => enable_passthrough_case_1_y_net_x2,
    kernel_result_valid_bus_7_1 => enable_passthrough_case_1_y_net_x1,
    kernel_result_valid_bus_8_1 => enable_passthrough_case_1_y_net_x0,
    kernel_result_valid_bus_9_1 => enable_passthrough_case_1_y_net,
    pixel_group_offset_0_2 => delay_2_q_net,
    pixel_group_offset_0_3 => delay_4_q_net,
    pixel_group_offset_0_4 => delay_6_q_net,
    pixel_group_offset_0_5 => delay_8_q_net,
    pixel_group_offset_0_6 => delay_10_q_net,
    pixel_group_offset_0_7 => delay_12_q_net,
    pixel_group_offset_0_8 => delay_14_q_net,
    pixel_group_offset_0_9 => delay_23_q_net,
    pixel_group_offset_0_10 => delay_16_q_net,
    pixel_group_offset_0_11 => delay_18_q_net,
    pixel_group_offset_0_12 => delay_20_q_net,
    pixel_group_offset_1_2 => delay_36_q_net,
    pixel_group_offset_1_3 => delay_42_q_net,
    pixel_group_offset_1_4 => delay_44_q_net,
    pixel_group_offset_1_5 => delay_46_q_net,
    pixel_group_offset_1_6 => delay_26_q_net,
    pixel_group_offset_1_7 => delay_28_q_net,
    pixel_group_offset_1_8 => delay_30_q_net,
    pixel_group_offset_1_9 => delay_39_q_net,
    pixel_group_offset_1_10 => delay_32_q_net,
    pixel_group_offset_1_11 => delay_34_q_net,
    pixel_group_offset_1_12 => delay_37_q_net,
    pixel_group_offset_2_2 => delay_60_q_net,
    pixel_group_offset_2_3 => delay_66_q_net,
    pixel_group_offset_2_4 => delay_68_q_net,
    pixel_group_offset_2_5 => delay_70_q_net,
    pixel_group_offset_2_6 => delay_50_q_net,
    pixel_group_offset_2_7 => delay_52_q_net,
    pixel_group_offset_2_8 => delay_54_q_net,
    pixel_group_offset_2_9 => delay_63_q_net,
    pixel_group_offset_2_10 => delay_56_q_net,
    pixel_group_offset_2_11 => delay_58_q_net,
    pixel_group_offset_2_12 => delay_61_q_net,
    pixel_group_offset_3_2 => delay_84_q_net,
    pixel_group_offset_3_3 => delay_90_q_net,
    pixel_group_offset_3_4 => delay_92_q_net,
    pixel_group_offset_3_5 => delay_94_q_net,
    pixel_group_offset_3_6 => delay_74_q_net,
    pixel_group_offset_3_7 => delay_76_q_net,
    pixel_group_offset_3_8 => delay_78_q_net,
    pixel_group_offset_3_9 => delay_87_q_net,
    pixel_group_offset_3_10 => delay_80_q_net,
    pixel_group_offset_3_11 => delay_82_q_net,
    pixel_group_offset_3_12 => delay_85_q_net,
    pixel_group_offset_4_2 => delay_108_q_net,
    pixel_group_offset_4_3 => delay_114_q_net,
    pixel_group_offset_4_4 => delay_116_q_net,
    pixel_group_offset_4_5 => delay_118_q_net,
    pixel_group_offset_4_6 => delay_98_q_net,
    pixel_group_offset_4_7 => delay_100_q_net,
    pixel_group_offset_4_8 => delay_102_q_net,
    pixel_group_offset_4_9 => delay_111_q_net,
    pixel_group_offset_4_10 => delay_104_q_net,
    pixel_group_offset_4_11 => delay_106_q_net,
    pixel_group_offset_4_12 => delay_109_q_net,
    weights_2 => delay_3_q_net,
    weights_3 => delay_5_q_net,
    weights_4 => delay_7_q_net,
    weights_5 => delay_9_q_net,
    weights_6 => delay_11_q_net,
    weights_7 => delay_13_q_net,
    weights_8 => delay_15_q_net,
    weights_9 => delay_24_q_net,
    weights_10 => delay_17_q_net,
    weights_11 => delay_19_q_net,
    weights_12 => delay_21_q_net,
    weights_13 => delay_25_q_net,
    weights_14 => delay_41_q_net,
    weights_15 => delay_43_q_net,
    weights_16 => delay_45_q_net,
    weights_17 => delay_47_q_net,
    weights_18 => delay_27_q_net,
    weights_19 => delay_29_q_net,
    weights_20 => delay_31_q_net,
    weights_21 => delay_40_q_net,
    weights_22 => delay_33_q_net,
    weights_23 => delay_35_q_net,
    weights_24 => delay_38_q_net,
    weights_25 => delay_49_q_net,
    weights_26 => delay_65_q_net,
    weights_27 => delay_67_q_net,
    weights_28 => delay_69_q_net,
    weights_29 => delay_71_q_net,
    weights_30 => delay_51_q_net,
    weights_31 => delay_53_q_net,
    weights_32 => delay_55_q_net,
    weights_33 => delay_64_q_net,
    weights_34 => delay_57_q_net,
    weights_35 => delay_59_q_net,
    weights_36 => delay_62_q_net,
    weights_37 => delay_73_q_net,
    weights_38 => delay_89_q_net,
    weights_39 => delay_91_q_net,
    weights_40 => delay_93_q_net,
    weights_41 => delay_95_q_net,
    weights_42 => delay_75_q_net,
    weights_43 => delay_77_q_net,
    weights_44 => delay_79_q_net,
    weights_45 => delay_88_q_net,
    weights_46 => delay_81_q_net,
    weights_47 => delay_83_q_net,
    weights_48 => delay_86_q_net,
    weights_49 => delay_97_q_net,
    weights_50 => delay_113_q_net,
    weights_51 => delay_115_q_net,
    weights_52 => delay_117_q_net,
    weights_53 => delay_119_q_net,
    weights_54 => delay_99_q_net,
    weights_55 => delay_101_q_net,
    weights_56 => delay_103_q_net,
    weights_57 => delay_112_q_net,
    weights_58 => delay_105_q_net,
    weights_59 => delay_107_q_net,
    weights_60 => delay_110_q_net,
    weights_61 => last_out_q_net,
    kernel_result_valid_bus_0_2 => enable_passthrough_case_0_y_net_x7,
    kernel_result_valid_bus_0_3 => enable_passthrough_case_0_y_net_x7,
    kernel_result_valid_bus_0_4 => enable_passthrough_case_0_y_net_x7,
    kernel_result_valid_bus_0_5 => enable_passthrough_case_0_y_net_x7,
    kernel_result_valid_bus_1_2 => enable_passthrough_case_0_y_net_x6,
    kernel_result_valid_bus_1_3 => enable_passthrough_case_0_y_net_x6,
    kernel_result_valid_bus_1_4 => enable_passthrough_case_0_y_net_x6,
    kernel_result_valid_bus_1_5 => enable_passthrough_case_1_y_net_x7,
    kernel_result_valid_bus_2_2 => enable_passthrough_case_0_y_net_x5,
    kernel_result_valid_bus_2_3 => enable_passthrough_case_0_y_net_x5,
    kernel_result_valid_bus_2_4 => enable_passthrough_case_1_y_net_x6,
    kernel_result_valid_bus_2_5 => enable_passthrough_case_1_y_net_x6,
    kernel_result_valid_bus_3_2 => enable_passthrough_case_0_y_net_x4,
    kernel_result_valid_bus_3_3 => enable_passthrough_case_1_y_net_x5,
    kernel_result_valid_bus_3_4 => enable_passthrough_case_1_y_net_x5,
    kernel_result_valid_bus_3_5 => enable_passthrough_case_1_y_net_x5,
    kernel_result_valid_bus_4_2 => enable_passthrough_case_1_y_net_x4,
    kernel_result_valid_bus_4_3 => enable_passthrough_case_1_y_net_x4,
    kernel_result_valid_bus_4_4 => enable_passthrough_case_1_y_net_x4,
    kernel_result_valid_bus_4_5 => enable_passthrough_case_1_y_net_x4,
    kernel_result_valid_bus_5_2 => enable_passthrough_case_1_y_net_x3,
    kernel_result_valid_bus_5_3 => enable_passthrough_case_1_y_net_x3,
    kernel_result_valid_bus_5_4 => enable_passthrough_case_1_y_net_x3,
    kernel_result_valid_bus_5_5 => enable_passthrough_case_1_y_net_x3,
    kernel_result_valid_bus_6_2 => enable_passthrough_case_1_y_net_x2,
    kernel_result_valid_bus_6_3 => enable_passthrough_case_1_y_net_x2,
    kernel_result_valid_bus_6_4 => enable_passthrough_case_1_y_net_x2,
    kernel_result_valid_bus_6_5 => enable_passthrough_case_0_y_net_x2,
    kernel_result_valid_bus_7_2 => enable_passthrough_case_1_y_net_x1,
    kernel_result_valid_bus_7_3 => enable_passthrough_case_1_y_net_x1,
    kernel_result_valid_bus_7_4 => enable_passthrough_case_0_y_net_x1,
    kernel_result_valid_bus_7_5 => enable_passthrough_case_0_y_net_x1,
    kernel_result_valid_bus_8_2 => enable_passthrough_case_1_y_net_x0,
    kernel_result_valid_bus_8_3 => enable_passthrough_case_0_y_net_x0,
    kernel_result_valid_bus_8_4 => enable_passthrough_case_0_y_net_x0,
    kernel_result_valid_bus_8_5 => enable_passthrough_case_0_y_net_x0,
    kernel_result_valid_bus_9_2 => enable_passthrough_case_0_y_net,
    kernel_result_valid_bus_9_3 => enable_passthrough_case_0_y_net,
    kernel_result_valid_bus_9_4 => enable_passthrough_case_0_y_net,
    kernel_result_valid_bus_9_5 => enable_passthrough_case_0_y_net
  );
  kernel_result_0 : entity xil_defaultlib.mh_kernel_result_0 
  port map (
    pixel_bus_input_offset_0_1 => delay_0_q_net,
    pixel_bus_input_offset_1_1 => delay_22_q_net,
    pixel_bus_input_offset_2_1 => delay_48_q_net,
    pixel_bus_input_offset_3_1 => delay_72_q_net,
    pixel_bus_input_offset_4_1 => delay_96_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_0_y_net_x7,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_2_q_net,
    pixel_bus_input_offset_0_3 => delay_4_q_net,
    pixel_bus_input_offset_0_4 => delay_6_q_net,
    pixel_bus_input_offset_0_5 => delay_8_q_net,
    pixel_bus_input_offset_0_6 => delay_10_q_net,
    pixel_bus_input_offset_0_7 => delay_12_q_net,
    pixel_bus_input_offset_0_8 => delay_14_q_net,
    pixel_bus_input_offset_0_9 => delay_23_q_net,
    pixel_bus_input_offset_0_10 => delay_16_q_net,
    pixel_bus_input_offset_0_11 => delay_18_q_net,
    pixel_bus_input_offset_0_12 => delay_20_q_net,
    pixel_bus_input_offset_1_2 => delay_36_q_net,
    pixel_bus_input_offset_1_3 => delay_42_q_net,
    pixel_bus_input_offset_1_4 => delay_44_q_net,
    pixel_bus_input_offset_1_5 => delay_46_q_net,
    pixel_bus_input_offset_1_6 => delay_26_q_net,
    pixel_bus_input_offset_1_7 => delay_28_q_net,
    pixel_bus_input_offset_1_8 => delay_30_q_net,
    pixel_bus_input_offset_1_9 => delay_39_q_net,
    pixel_bus_input_offset_1_10 => delay_32_q_net,
    pixel_bus_input_offset_1_11 => delay_34_q_net,
    pixel_bus_input_offset_1_12 => delay_37_q_net,
    pixel_bus_input_offset_2_2 => delay_60_q_net,
    pixel_bus_input_offset_2_3 => delay_66_q_net,
    pixel_bus_input_offset_2_4 => delay_68_q_net,
    pixel_bus_input_offset_2_5 => delay_70_q_net,
    pixel_bus_input_offset_2_6 => delay_50_q_net,
    pixel_bus_input_offset_2_7 => delay_52_q_net,
    pixel_bus_input_offset_2_8 => delay_54_q_net,
    pixel_bus_input_offset_2_9 => delay_63_q_net,
    pixel_bus_input_offset_2_10 => delay_56_q_net,
    pixel_bus_input_offset_2_11 => delay_58_q_net,
    pixel_bus_input_offset_2_12 => delay_61_q_net,
    pixel_bus_input_offset_3_2 => delay_84_q_net,
    pixel_bus_input_offset_3_3 => delay_90_q_net,
    pixel_bus_input_offset_3_4 => delay_92_q_net,
    pixel_bus_input_offset_3_5 => delay_94_q_net,
    pixel_bus_input_offset_3_6 => delay_74_q_net,
    pixel_bus_input_offset_3_7 => delay_76_q_net,
    pixel_bus_input_offset_3_8 => delay_78_q_net,
    pixel_bus_input_offset_3_9 => delay_87_q_net,
    pixel_bus_input_offset_3_10 => delay_80_q_net,
    pixel_bus_input_offset_3_11 => delay_82_q_net,
    pixel_bus_input_offset_3_12 => delay_85_q_net,
    pixel_bus_input_offset_4_2 => delay_108_q_net,
    pixel_bus_input_offset_4_3 => delay_114_q_net,
    pixel_bus_input_offset_4_4 => delay_116_q_net,
    pixel_bus_input_offset_4_5 => delay_118_q_net,
    pixel_bus_input_offset_4_6 => delay_98_q_net,
    pixel_bus_input_offset_4_7 => delay_100_q_net,
    pixel_bus_input_offset_4_8 => delay_102_q_net,
    pixel_bus_input_offset_4_9 => delay_111_q_net,
    pixel_bus_input_offset_4_10 => delay_104_q_net,
    pixel_bus_input_offset_4_11 => delay_106_q_net,
    pixel_bus_input_offset_4_12 => delay_109_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x6,
    valid_kernel_output => delay_enable_4_q_net_x5
  );
  kernel_result_1 : entity xil_defaultlib.mh_kernel_result_1 
  port map (
    pixel_bus_input_offset_0_1 => delay_22_q_net,
    pixel_bus_input_offset_1_1 => delay_48_q_net,
    pixel_bus_input_offset_2_1 => delay_72_q_net,
    pixel_bus_input_offset_3_1 => delay_96_q_net,
    pixel_bus_input_offset_4_1 => delay_0_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_0_y_net_x6,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_36_q_net,
    pixel_bus_input_offset_0_3 => delay_42_q_net,
    pixel_bus_input_offset_0_4 => delay_44_q_net,
    pixel_bus_input_offset_0_5 => delay_46_q_net,
    pixel_bus_input_offset_0_6 => delay_26_q_net,
    pixel_bus_input_offset_0_7 => delay_28_q_net,
    pixel_bus_input_offset_0_8 => delay_30_q_net,
    pixel_bus_input_offset_0_9 => delay_39_q_net,
    pixel_bus_input_offset_0_10 => delay_32_q_net,
    pixel_bus_input_offset_0_11 => delay_34_q_net,
    pixel_bus_input_offset_0_12 => delay_37_q_net,
    pixel_bus_input_offset_1_2 => delay_60_q_net,
    pixel_bus_input_offset_1_3 => delay_66_q_net,
    pixel_bus_input_offset_1_4 => delay_68_q_net,
    pixel_bus_input_offset_1_5 => delay_70_q_net,
    pixel_bus_input_offset_1_6 => delay_50_q_net,
    pixel_bus_input_offset_1_7 => delay_52_q_net,
    pixel_bus_input_offset_1_8 => delay_54_q_net,
    pixel_bus_input_offset_1_9 => delay_63_q_net,
    pixel_bus_input_offset_1_10 => delay_56_q_net,
    pixel_bus_input_offset_1_11 => delay_58_q_net,
    pixel_bus_input_offset_1_12 => delay_61_q_net,
    pixel_bus_input_offset_2_2 => delay_84_q_net,
    pixel_bus_input_offset_2_3 => delay_90_q_net,
    pixel_bus_input_offset_2_4 => delay_92_q_net,
    pixel_bus_input_offset_2_5 => delay_94_q_net,
    pixel_bus_input_offset_2_6 => delay_74_q_net,
    pixel_bus_input_offset_2_7 => delay_76_q_net,
    pixel_bus_input_offset_2_8 => delay_78_q_net,
    pixel_bus_input_offset_2_9 => delay_87_q_net,
    pixel_bus_input_offset_2_10 => delay_80_q_net,
    pixel_bus_input_offset_2_11 => delay_82_q_net,
    pixel_bus_input_offset_2_12 => delay_85_q_net,
    pixel_bus_input_offset_3_2 => delay_108_q_net,
    pixel_bus_input_offset_3_3 => delay_114_q_net,
    pixel_bus_input_offset_3_4 => delay_116_q_net,
    pixel_bus_input_offset_3_5 => delay_118_q_net,
    pixel_bus_input_offset_3_6 => delay_98_q_net,
    pixel_bus_input_offset_3_7 => delay_100_q_net,
    pixel_bus_input_offset_3_8 => delay_102_q_net,
    pixel_bus_input_offset_3_9 => delay_111_q_net,
    pixel_bus_input_offset_3_10 => delay_104_q_net,
    pixel_bus_input_offset_3_11 => delay_106_q_net,
    pixel_bus_input_offset_3_12 => delay_109_q_net,
    pixel_bus_input_offset_4_2 => delay_2_q_net,
    pixel_bus_input_offset_4_3 => delay_4_q_net,
    pixel_bus_input_offset_4_4 => delay_6_q_net,
    pixel_bus_input_offset_4_5 => delay_8_q_net,
    pixel_bus_input_offset_4_6 => delay_10_q_net,
    pixel_bus_input_offset_4_7 => delay_12_q_net,
    pixel_bus_input_offset_4_8 => delay_14_q_net,
    pixel_bus_input_offset_4_9 => delay_23_q_net,
    pixel_bus_input_offset_4_10 => delay_16_q_net,
    pixel_bus_input_offset_4_11 => delay_18_q_net,
    pixel_bus_input_offset_4_12 => delay_20_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_5 => enable_passthrough_case_1_y_net_x7,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x5,
    valid_kernel_output => delay_enable_4_q_net_x4
  );
  kernel_result_2 : entity xil_defaultlib.mh_kernel_result_2 
  port map (
    pixel_bus_input_offset_0_1 => delay_48_q_net,
    pixel_bus_input_offset_1_1 => delay_72_q_net,
    pixel_bus_input_offset_2_1 => delay_96_q_net,
    pixel_bus_input_offset_3_1 => delay_0_q_net,
    pixel_bus_input_offset_4_1 => delay_22_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_0_y_net_x5,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_60_q_net,
    pixel_bus_input_offset_0_3 => delay_66_q_net,
    pixel_bus_input_offset_0_4 => delay_68_q_net,
    pixel_bus_input_offset_0_5 => delay_70_q_net,
    pixel_bus_input_offset_0_6 => delay_50_q_net,
    pixel_bus_input_offset_0_7 => delay_52_q_net,
    pixel_bus_input_offset_0_8 => delay_54_q_net,
    pixel_bus_input_offset_0_9 => delay_63_q_net,
    pixel_bus_input_offset_0_10 => delay_56_q_net,
    pixel_bus_input_offset_0_11 => delay_58_q_net,
    pixel_bus_input_offset_0_12 => delay_61_q_net,
    pixel_bus_input_offset_1_2 => delay_84_q_net,
    pixel_bus_input_offset_1_3 => delay_90_q_net,
    pixel_bus_input_offset_1_4 => delay_92_q_net,
    pixel_bus_input_offset_1_5 => delay_94_q_net,
    pixel_bus_input_offset_1_6 => delay_74_q_net,
    pixel_bus_input_offset_1_7 => delay_76_q_net,
    pixel_bus_input_offset_1_8 => delay_78_q_net,
    pixel_bus_input_offset_1_9 => delay_87_q_net,
    pixel_bus_input_offset_1_10 => delay_80_q_net,
    pixel_bus_input_offset_1_11 => delay_82_q_net,
    pixel_bus_input_offset_1_12 => delay_85_q_net,
    pixel_bus_input_offset_2_2 => delay_108_q_net,
    pixel_bus_input_offset_2_3 => delay_114_q_net,
    pixel_bus_input_offset_2_4 => delay_116_q_net,
    pixel_bus_input_offset_2_5 => delay_118_q_net,
    pixel_bus_input_offset_2_6 => delay_98_q_net,
    pixel_bus_input_offset_2_7 => delay_100_q_net,
    pixel_bus_input_offset_2_8 => delay_102_q_net,
    pixel_bus_input_offset_2_9 => delay_111_q_net,
    pixel_bus_input_offset_2_10 => delay_104_q_net,
    pixel_bus_input_offset_2_11 => delay_106_q_net,
    pixel_bus_input_offset_2_12 => delay_109_q_net,
    pixel_bus_input_offset_3_2 => delay_2_q_net,
    pixel_bus_input_offset_3_3 => delay_4_q_net,
    pixel_bus_input_offset_3_4 => delay_6_q_net,
    pixel_bus_input_offset_3_5 => delay_8_q_net,
    pixel_bus_input_offset_3_6 => delay_10_q_net,
    pixel_bus_input_offset_3_7 => delay_12_q_net,
    pixel_bus_input_offset_3_8 => delay_14_q_net,
    pixel_bus_input_offset_3_9 => delay_23_q_net,
    pixel_bus_input_offset_3_10 => delay_16_q_net,
    pixel_bus_input_offset_3_11 => delay_18_q_net,
    pixel_bus_input_offset_3_12 => delay_20_q_net,
    pixel_bus_input_offset_4_2 => delay_36_q_net,
    pixel_bus_input_offset_4_3 => delay_42_q_net,
    pixel_bus_input_offset_4_4 => delay_44_q_net,
    pixel_bus_input_offset_4_5 => delay_46_q_net,
    pixel_bus_input_offset_4_6 => delay_26_q_net,
    pixel_bus_input_offset_4_7 => delay_28_q_net,
    pixel_bus_input_offset_4_8 => delay_30_q_net,
    pixel_bus_input_offset_4_9 => delay_39_q_net,
    pixel_bus_input_offset_4_10 => delay_32_q_net,
    pixel_bus_input_offset_4_11 => delay_34_q_net,
    pixel_bus_input_offset_4_12 => delay_37_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_4 => enable_passthrough_case_1_y_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x4,
    valid_kernel_output => delay_enable_4_q_net_x3
  );
  kernel_result_3 : entity xil_defaultlib.mh_kernel_result_3 
  port map (
    pixel_bus_input_offset_0_1 => delay_72_q_net,
    pixel_bus_input_offset_1_1 => delay_96_q_net,
    pixel_bus_input_offset_2_1 => delay_0_q_net,
    pixel_bus_input_offset_3_1 => delay_22_q_net,
    pixel_bus_input_offset_4_1 => delay_48_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_0_y_net_x4,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_84_q_net,
    pixel_bus_input_offset_0_3 => delay_90_q_net,
    pixel_bus_input_offset_0_4 => delay_92_q_net,
    pixel_bus_input_offset_0_5 => delay_94_q_net,
    pixel_bus_input_offset_0_6 => delay_74_q_net,
    pixel_bus_input_offset_0_7 => delay_76_q_net,
    pixel_bus_input_offset_0_8 => delay_78_q_net,
    pixel_bus_input_offset_0_9 => delay_87_q_net,
    pixel_bus_input_offset_0_10 => delay_80_q_net,
    pixel_bus_input_offset_0_11 => delay_82_q_net,
    pixel_bus_input_offset_0_12 => delay_85_q_net,
    pixel_bus_input_offset_1_2 => delay_108_q_net,
    pixel_bus_input_offset_1_3 => delay_114_q_net,
    pixel_bus_input_offset_1_4 => delay_116_q_net,
    pixel_bus_input_offset_1_5 => delay_118_q_net,
    pixel_bus_input_offset_1_6 => delay_98_q_net,
    pixel_bus_input_offset_1_7 => delay_100_q_net,
    pixel_bus_input_offset_1_8 => delay_102_q_net,
    pixel_bus_input_offset_1_9 => delay_111_q_net,
    pixel_bus_input_offset_1_10 => delay_104_q_net,
    pixel_bus_input_offset_1_11 => delay_106_q_net,
    pixel_bus_input_offset_1_12 => delay_109_q_net,
    pixel_bus_input_offset_2_2 => delay_2_q_net,
    pixel_bus_input_offset_2_3 => delay_4_q_net,
    pixel_bus_input_offset_2_4 => delay_6_q_net,
    pixel_bus_input_offset_2_5 => delay_8_q_net,
    pixel_bus_input_offset_2_6 => delay_10_q_net,
    pixel_bus_input_offset_2_7 => delay_12_q_net,
    pixel_bus_input_offset_2_8 => delay_14_q_net,
    pixel_bus_input_offset_2_9 => delay_23_q_net,
    pixel_bus_input_offset_2_10 => delay_16_q_net,
    pixel_bus_input_offset_2_11 => delay_18_q_net,
    pixel_bus_input_offset_2_12 => delay_20_q_net,
    pixel_bus_input_offset_3_2 => delay_36_q_net,
    pixel_bus_input_offset_3_3 => delay_42_q_net,
    pixel_bus_input_offset_3_4 => delay_44_q_net,
    pixel_bus_input_offset_3_5 => delay_46_q_net,
    pixel_bus_input_offset_3_6 => delay_26_q_net,
    pixel_bus_input_offset_3_7 => delay_28_q_net,
    pixel_bus_input_offset_3_8 => delay_30_q_net,
    pixel_bus_input_offset_3_9 => delay_39_q_net,
    pixel_bus_input_offset_3_10 => delay_32_q_net,
    pixel_bus_input_offset_3_11 => delay_34_q_net,
    pixel_bus_input_offset_3_12 => delay_37_q_net,
    pixel_bus_input_offset_4_2 => delay_60_q_net,
    pixel_bus_input_offset_4_3 => delay_66_q_net,
    pixel_bus_input_offset_4_4 => delay_68_q_net,
    pixel_bus_input_offset_4_5 => delay_70_q_net,
    pixel_bus_input_offset_4_6 => delay_50_q_net,
    pixel_bus_input_offset_4_7 => delay_52_q_net,
    pixel_bus_input_offset_4_8 => delay_54_q_net,
    pixel_bus_input_offset_4_9 => delay_63_q_net,
    pixel_bus_input_offset_4_10 => delay_56_q_net,
    pixel_bus_input_offset_4_11 => delay_58_q_net,
    pixel_bus_input_offset_4_12 => delay_61_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_3 => enable_passthrough_case_1_y_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x3,
    valid_kernel_output => delay_enable_4_q_net_x2
  );
  kernel_result_4 : entity xil_defaultlib.mh_kernel_result_4 
  port map (
    pixel_bus_input_offset_0_1 => delay_96_q_net,
    pixel_bus_input_offset_1_1 => delay_0_q_net,
    pixel_bus_input_offset_2_1 => delay_22_q_net,
    pixel_bus_input_offset_3_1 => delay_48_q_net,
    pixel_bus_input_offset_4_1 => delay_72_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_0_y_net_x3,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_108_q_net,
    pixel_bus_input_offset_0_3 => delay_114_q_net,
    pixel_bus_input_offset_0_4 => delay_116_q_net,
    pixel_bus_input_offset_0_5 => delay_118_q_net,
    pixel_bus_input_offset_0_6 => delay_98_q_net,
    pixel_bus_input_offset_0_7 => delay_100_q_net,
    pixel_bus_input_offset_0_8 => delay_102_q_net,
    pixel_bus_input_offset_0_9 => delay_111_q_net,
    pixel_bus_input_offset_0_10 => delay_104_q_net,
    pixel_bus_input_offset_0_11 => delay_106_q_net,
    pixel_bus_input_offset_0_12 => delay_109_q_net,
    pixel_bus_input_offset_1_2 => delay_2_q_net,
    pixel_bus_input_offset_1_3 => delay_4_q_net,
    pixel_bus_input_offset_1_4 => delay_6_q_net,
    pixel_bus_input_offset_1_5 => delay_8_q_net,
    pixel_bus_input_offset_1_6 => delay_10_q_net,
    pixel_bus_input_offset_1_7 => delay_12_q_net,
    pixel_bus_input_offset_1_8 => delay_14_q_net,
    pixel_bus_input_offset_1_9 => delay_23_q_net,
    pixel_bus_input_offset_1_10 => delay_16_q_net,
    pixel_bus_input_offset_1_11 => delay_18_q_net,
    pixel_bus_input_offset_1_12 => delay_20_q_net,
    pixel_bus_input_offset_2_2 => delay_36_q_net,
    pixel_bus_input_offset_2_3 => delay_42_q_net,
    pixel_bus_input_offset_2_4 => delay_44_q_net,
    pixel_bus_input_offset_2_5 => delay_46_q_net,
    pixel_bus_input_offset_2_6 => delay_26_q_net,
    pixel_bus_input_offset_2_7 => delay_28_q_net,
    pixel_bus_input_offset_2_8 => delay_30_q_net,
    pixel_bus_input_offset_2_9 => delay_39_q_net,
    pixel_bus_input_offset_2_10 => delay_32_q_net,
    pixel_bus_input_offset_2_11 => delay_34_q_net,
    pixel_bus_input_offset_2_12 => delay_37_q_net,
    pixel_bus_input_offset_3_2 => delay_60_q_net,
    pixel_bus_input_offset_3_3 => delay_66_q_net,
    pixel_bus_input_offset_3_4 => delay_68_q_net,
    pixel_bus_input_offset_3_5 => delay_70_q_net,
    pixel_bus_input_offset_3_6 => delay_50_q_net,
    pixel_bus_input_offset_3_7 => delay_52_q_net,
    pixel_bus_input_offset_3_8 => delay_54_q_net,
    pixel_bus_input_offset_3_9 => delay_63_q_net,
    pixel_bus_input_offset_3_10 => delay_56_q_net,
    pixel_bus_input_offset_3_11 => delay_58_q_net,
    pixel_bus_input_offset_3_12 => delay_61_q_net,
    pixel_bus_input_offset_4_2 => delay_84_q_net,
    pixel_bus_input_offset_4_3 => delay_90_q_net,
    pixel_bus_input_offset_4_4 => delay_92_q_net,
    pixel_bus_input_offset_4_5 => delay_94_q_net,
    pixel_bus_input_offset_4_6 => delay_74_q_net,
    pixel_bus_input_offset_4_7 => delay_76_q_net,
    pixel_bus_input_offset_4_8 => delay_78_q_net,
    pixel_bus_input_offset_4_9 => delay_87_q_net,
    pixel_bus_input_offset_4_10 => delay_80_q_net,
    pixel_bus_input_offset_4_11 => delay_82_q_net,
    pixel_bus_input_offset_4_12 => delay_85_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_2 => enable_passthrough_case_1_y_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x2,
    valid_kernel_output => delay_enable_4_q_net_x1
  );
  kernel_result_5 : entity xil_defaultlib.mh_kernel_result_5 
  port map (
    pixel_bus_input_offset_0_1 => delay_0_q_net,
    pixel_bus_input_offset_1_1 => delay_22_q_net,
    pixel_bus_input_offset_2_1 => delay_48_q_net,
    pixel_bus_input_offset_3_1 => delay_72_q_net,
    pixel_bus_input_offset_4_1 => delay_96_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_1_y_net_x3,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_2_q_net,
    pixel_bus_input_offset_0_3 => delay_4_q_net,
    pixel_bus_input_offset_0_4 => delay_6_q_net,
    pixel_bus_input_offset_0_5 => delay_8_q_net,
    pixel_bus_input_offset_0_6 => delay_10_q_net,
    pixel_bus_input_offset_0_7 => delay_12_q_net,
    pixel_bus_input_offset_0_8 => delay_14_q_net,
    pixel_bus_input_offset_0_9 => delay_23_q_net,
    pixel_bus_input_offset_0_10 => delay_16_q_net,
    pixel_bus_input_offset_0_11 => delay_18_q_net,
    pixel_bus_input_offset_0_12 => delay_20_q_net,
    pixel_bus_input_offset_1_2 => delay_36_q_net,
    pixel_bus_input_offset_1_3 => delay_42_q_net,
    pixel_bus_input_offset_1_4 => delay_44_q_net,
    pixel_bus_input_offset_1_5 => delay_46_q_net,
    pixel_bus_input_offset_1_6 => delay_26_q_net,
    pixel_bus_input_offset_1_7 => delay_28_q_net,
    pixel_bus_input_offset_1_8 => delay_30_q_net,
    pixel_bus_input_offset_1_9 => delay_39_q_net,
    pixel_bus_input_offset_1_10 => delay_32_q_net,
    pixel_bus_input_offset_1_11 => delay_34_q_net,
    pixel_bus_input_offset_1_12 => delay_37_q_net,
    pixel_bus_input_offset_2_2 => delay_60_q_net,
    pixel_bus_input_offset_2_3 => delay_66_q_net,
    pixel_bus_input_offset_2_4 => delay_68_q_net,
    pixel_bus_input_offset_2_5 => delay_70_q_net,
    pixel_bus_input_offset_2_6 => delay_50_q_net,
    pixel_bus_input_offset_2_7 => delay_52_q_net,
    pixel_bus_input_offset_2_8 => delay_54_q_net,
    pixel_bus_input_offset_2_9 => delay_63_q_net,
    pixel_bus_input_offset_2_10 => delay_56_q_net,
    pixel_bus_input_offset_2_11 => delay_58_q_net,
    pixel_bus_input_offset_2_12 => delay_61_q_net,
    pixel_bus_input_offset_3_2 => delay_84_q_net,
    pixel_bus_input_offset_3_3 => delay_90_q_net,
    pixel_bus_input_offset_3_4 => delay_92_q_net,
    pixel_bus_input_offset_3_5 => delay_94_q_net,
    pixel_bus_input_offset_3_6 => delay_74_q_net,
    pixel_bus_input_offset_3_7 => delay_76_q_net,
    pixel_bus_input_offset_3_8 => delay_78_q_net,
    pixel_bus_input_offset_3_9 => delay_87_q_net,
    pixel_bus_input_offset_3_10 => delay_80_q_net,
    pixel_bus_input_offset_3_11 => delay_82_q_net,
    pixel_bus_input_offset_3_12 => delay_85_q_net,
    pixel_bus_input_offset_4_2 => delay_108_q_net,
    pixel_bus_input_offset_4_3 => delay_114_q_net,
    pixel_bus_input_offset_4_4 => delay_116_q_net,
    pixel_bus_input_offset_4_5 => delay_118_q_net,
    pixel_bus_input_offset_4_6 => delay_98_q_net,
    pixel_bus_input_offset_4_7 => delay_100_q_net,
    pixel_bus_input_offset_4_8 => delay_102_q_net,
    pixel_bus_input_offset_4_9 => delay_111_q_net,
    pixel_bus_input_offset_4_10 => delay_104_q_net,
    pixel_bus_input_offset_4_11 => delay_106_q_net,
    pixel_bus_input_offset_4_12 => delay_109_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x1,
    valid_kernel_output => delay_enable_4_q_net_x0
  );
  kernel_result_6 : entity xil_defaultlib.mh_kernel_result_6 
  port map (
    pixel_bus_input_offset_0_1 => delay_22_q_net,
    pixel_bus_input_offset_1_1 => delay_48_q_net,
    pixel_bus_input_offset_2_1 => delay_72_q_net,
    pixel_bus_input_offset_3_1 => delay_96_q_net,
    pixel_bus_input_offset_4_1 => delay_0_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_1_y_net_x2,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_36_q_net,
    pixel_bus_input_offset_0_3 => delay_42_q_net,
    pixel_bus_input_offset_0_4 => delay_44_q_net,
    pixel_bus_input_offset_0_5 => delay_46_q_net,
    pixel_bus_input_offset_0_6 => delay_26_q_net,
    pixel_bus_input_offset_0_7 => delay_28_q_net,
    pixel_bus_input_offset_0_8 => delay_30_q_net,
    pixel_bus_input_offset_0_9 => delay_39_q_net,
    pixel_bus_input_offset_0_10 => delay_32_q_net,
    pixel_bus_input_offset_0_11 => delay_34_q_net,
    pixel_bus_input_offset_0_12 => delay_37_q_net,
    pixel_bus_input_offset_1_2 => delay_60_q_net,
    pixel_bus_input_offset_1_3 => delay_66_q_net,
    pixel_bus_input_offset_1_4 => delay_68_q_net,
    pixel_bus_input_offset_1_5 => delay_70_q_net,
    pixel_bus_input_offset_1_6 => delay_50_q_net,
    pixel_bus_input_offset_1_7 => delay_52_q_net,
    pixel_bus_input_offset_1_8 => delay_54_q_net,
    pixel_bus_input_offset_1_9 => delay_63_q_net,
    pixel_bus_input_offset_1_10 => delay_56_q_net,
    pixel_bus_input_offset_1_11 => delay_58_q_net,
    pixel_bus_input_offset_1_12 => delay_61_q_net,
    pixel_bus_input_offset_2_2 => delay_84_q_net,
    pixel_bus_input_offset_2_3 => delay_90_q_net,
    pixel_bus_input_offset_2_4 => delay_92_q_net,
    pixel_bus_input_offset_2_5 => delay_94_q_net,
    pixel_bus_input_offset_2_6 => delay_74_q_net,
    pixel_bus_input_offset_2_7 => delay_76_q_net,
    pixel_bus_input_offset_2_8 => delay_78_q_net,
    pixel_bus_input_offset_2_9 => delay_87_q_net,
    pixel_bus_input_offset_2_10 => delay_80_q_net,
    pixel_bus_input_offset_2_11 => delay_82_q_net,
    pixel_bus_input_offset_2_12 => delay_85_q_net,
    pixel_bus_input_offset_3_2 => delay_108_q_net,
    pixel_bus_input_offset_3_3 => delay_114_q_net,
    pixel_bus_input_offset_3_4 => delay_116_q_net,
    pixel_bus_input_offset_3_5 => delay_118_q_net,
    pixel_bus_input_offset_3_6 => delay_98_q_net,
    pixel_bus_input_offset_3_7 => delay_100_q_net,
    pixel_bus_input_offset_3_8 => delay_102_q_net,
    pixel_bus_input_offset_3_9 => delay_111_q_net,
    pixel_bus_input_offset_3_10 => delay_104_q_net,
    pixel_bus_input_offset_3_11 => delay_106_q_net,
    pixel_bus_input_offset_3_12 => delay_109_q_net,
    pixel_bus_input_offset_4_2 => delay_2_q_net,
    pixel_bus_input_offset_4_3 => delay_4_q_net,
    pixel_bus_input_offset_4_4 => delay_6_q_net,
    pixel_bus_input_offset_4_5 => delay_8_q_net,
    pixel_bus_input_offset_4_6 => delay_10_q_net,
    pixel_bus_input_offset_4_7 => delay_12_q_net,
    pixel_bus_input_offset_4_8 => delay_14_q_net,
    pixel_bus_input_offset_4_9 => delay_23_q_net,
    pixel_bus_input_offset_4_10 => delay_16_q_net,
    pixel_bus_input_offset_4_11 => delay_18_q_net,
    pixel_bus_input_offset_4_12 => delay_20_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_5 => enable_passthrough_case_0_y_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x0,
    valid_kernel_output => delay_enable_4_q_net
  );
  kernel_result_7 : entity xil_defaultlib.mh_kernel_result_7 
  port map (
    pixel_bus_input_offset_0_1 => delay_48_q_net,
    pixel_bus_input_offset_1_1 => delay_72_q_net,
    pixel_bus_input_offset_2_1 => delay_96_q_net,
    pixel_bus_input_offset_3_1 => delay_0_q_net,
    pixel_bus_input_offset_4_1 => delay_22_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_1_y_net_x1,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_60_q_net,
    pixel_bus_input_offset_0_3 => delay_66_q_net,
    pixel_bus_input_offset_0_4 => delay_68_q_net,
    pixel_bus_input_offset_0_5 => delay_70_q_net,
    pixel_bus_input_offset_0_6 => delay_50_q_net,
    pixel_bus_input_offset_0_7 => delay_52_q_net,
    pixel_bus_input_offset_0_8 => delay_54_q_net,
    pixel_bus_input_offset_0_9 => delay_63_q_net,
    pixel_bus_input_offset_0_10 => delay_56_q_net,
    pixel_bus_input_offset_0_11 => delay_58_q_net,
    pixel_bus_input_offset_0_12 => delay_61_q_net,
    pixel_bus_input_offset_1_2 => delay_84_q_net,
    pixel_bus_input_offset_1_3 => delay_90_q_net,
    pixel_bus_input_offset_1_4 => delay_92_q_net,
    pixel_bus_input_offset_1_5 => delay_94_q_net,
    pixel_bus_input_offset_1_6 => delay_74_q_net,
    pixel_bus_input_offset_1_7 => delay_76_q_net,
    pixel_bus_input_offset_1_8 => delay_78_q_net,
    pixel_bus_input_offset_1_9 => delay_87_q_net,
    pixel_bus_input_offset_1_10 => delay_80_q_net,
    pixel_bus_input_offset_1_11 => delay_82_q_net,
    pixel_bus_input_offset_1_12 => delay_85_q_net,
    pixel_bus_input_offset_2_2 => delay_108_q_net,
    pixel_bus_input_offset_2_3 => delay_114_q_net,
    pixel_bus_input_offset_2_4 => delay_116_q_net,
    pixel_bus_input_offset_2_5 => delay_118_q_net,
    pixel_bus_input_offset_2_6 => delay_98_q_net,
    pixel_bus_input_offset_2_7 => delay_100_q_net,
    pixel_bus_input_offset_2_8 => delay_102_q_net,
    pixel_bus_input_offset_2_9 => delay_111_q_net,
    pixel_bus_input_offset_2_10 => delay_104_q_net,
    pixel_bus_input_offset_2_11 => delay_106_q_net,
    pixel_bus_input_offset_2_12 => delay_109_q_net,
    pixel_bus_input_offset_3_2 => delay_2_q_net,
    pixel_bus_input_offset_3_3 => delay_4_q_net,
    pixel_bus_input_offset_3_4 => delay_6_q_net,
    pixel_bus_input_offset_3_5 => delay_8_q_net,
    pixel_bus_input_offset_3_6 => delay_10_q_net,
    pixel_bus_input_offset_3_7 => delay_12_q_net,
    pixel_bus_input_offset_3_8 => delay_14_q_net,
    pixel_bus_input_offset_3_9 => delay_23_q_net,
    pixel_bus_input_offset_3_10 => delay_16_q_net,
    pixel_bus_input_offset_3_11 => delay_18_q_net,
    pixel_bus_input_offset_3_12 => delay_20_q_net,
    pixel_bus_input_offset_4_2 => delay_36_q_net,
    pixel_bus_input_offset_4_3 => delay_42_q_net,
    pixel_bus_input_offset_4_4 => delay_44_q_net,
    pixel_bus_input_offset_4_5 => delay_46_q_net,
    pixel_bus_input_offset_4_6 => delay_26_q_net,
    pixel_bus_input_offset_4_7 => delay_28_q_net,
    pixel_bus_input_offset_4_8 => delay_30_q_net,
    pixel_bus_input_offset_4_9 => delay_39_q_net,
    pixel_bus_input_offset_4_10 => delay_32_q_net,
    pixel_bus_input_offset_4_11 => delay_34_q_net,
    pixel_bus_input_offset_4_12 => delay_37_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_4 => enable_passthrough_case_0_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net,
    valid_kernel_output => delay_enable_4_q_net_x8
  );
  kernel_result_8 : entity xil_defaultlib.mh_kernel_result_8 
  port map (
    pixel_bus_input_offset_0_1 => delay_72_q_net,
    pixel_bus_input_offset_1_1 => delay_96_q_net,
    pixel_bus_input_offset_2_1 => delay_0_q_net,
    pixel_bus_input_offset_3_1 => delay_22_q_net,
    pixel_bus_input_offset_4_1 => delay_48_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_1_y_net_x0,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_84_q_net,
    pixel_bus_input_offset_0_3 => delay_90_q_net,
    pixel_bus_input_offset_0_4 => delay_92_q_net,
    pixel_bus_input_offset_0_5 => delay_94_q_net,
    pixel_bus_input_offset_0_6 => delay_74_q_net,
    pixel_bus_input_offset_0_7 => delay_76_q_net,
    pixel_bus_input_offset_0_8 => delay_78_q_net,
    pixel_bus_input_offset_0_9 => delay_87_q_net,
    pixel_bus_input_offset_0_10 => delay_80_q_net,
    pixel_bus_input_offset_0_11 => delay_82_q_net,
    pixel_bus_input_offset_0_12 => delay_85_q_net,
    pixel_bus_input_offset_1_2 => delay_108_q_net,
    pixel_bus_input_offset_1_3 => delay_114_q_net,
    pixel_bus_input_offset_1_4 => delay_116_q_net,
    pixel_bus_input_offset_1_5 => delay_118_q_net,
    pixel_bus_input_offset_1_6 => delay_98_q_net,
    pixel_bus_input_offset_1_7 => delay_100_q_net,
    pixel_bus_input_offset_1_8 => delay_102_q_net,
    pixel_bus_input_offset_1_9 => delay_111_q_net,
    pixel_bus_input_offset_1_10 => delay_104_q_net,
    pixel_bus_input_offset_1_11 => delay_106_q_net,
    pixel_bus_input_offset_1_12 => delay_109_q_net,
    pixel_bus_input_offset_2_2 => delay_2_q_net,
    pixel_bus_input_offset_2_3 => delay_4_q_net,
    pixel_bus_input_offset_2_4 => delay_6_q_net,
    pixel_bus_input_offset_2_5 => delay_8_q_net,
    pixel_bus_input_offset_2_6 => delay_10_q_net,
    pixel_bus_input_offset_2_7 => delay_12_q_net,
    pixel_bus_input_offset_2_8 => delay_14_q_net,
    pixel_bus_input_offset_2_9 => delay_23_q_net,
    pixel_bus_input_offset_2_10 => delay_16_q_net,
    pixel_bus_input_offset_2_11 => delay_18_q_net,
    pixel_bus_input_offset_2_12 => delay_20_q_net,
    pixel_bus_input_offset_3_2 => delay_36_q_net,
    pixel_bus_input_offset_3_3 => delay_42_q_net,
    pixel_bus_input_offset_3_4 => delay_44_q_net,
    pixel_bus_input_offset_3_5 => delay_46_q_net,
    pixel_bus_input_offset_3_6 => delay_26_q_net,
    pixel_bus_input_offset_3_7 => delay_28_q_net,
    pixel_bus_input_offset_3_8 => delay_30_q_net,
    pixel_bus_input_offset_3_9 => delay_39_q_net,
    pixel_bus_input_offset_3_10 => delay_32_q_net,
    pixel_bus_input_offset_3_11 => delay_34_q_net,
    pixel_bus_input_offset_3_12 => delay_37_q_net,
    pixel_bus_input_offset_4_2 => delay_60_q_net,
    pixel_bus_input_offset_4_3 => delay_66_q_net,
    pixel_bus_input_offset_4_4 => delay_68_q_net,
    pixel_bus_input_offset_4_5 => delay_70_q_net,
    pixel_bus_input_offset_4_6 => delay_50_q_net,
    pixel_bus_input_offset_4_7 => delay_52_q_net,
    pixel_bus_input_offset_4_8 => delay_54_q_net,
    pixel_bus_input_offset_4_9 => delay_63_q_net,
    pixel_bus_input_offset_4_10 => delay_56_q_net,
    pixel_bus_input_offset_4_11 => delay_58_q_net,
    pixel_bus_input_offset_4_12 => delay_61_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_3 => enable_passthrough_case_0_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x8,
    valid_kernel_output => delay_enable_4_q_net_x7
  );
  kernel_result_9 : entity xil_defaultlib.mh_kernel_result_9 
  port map (
    pixel_bus_input_offset_0_1 => delay_96_q_net,
    pixel_bus_input_offset_1_1 => delay_0_q_net,
    pixel_bus_input_offset_2_1 => delay_22_q_net,
    pixel_bus_input_offset_3_1 => delay_48_q_net,
    pixel_bus_input_offset_4_1 => delay_72_q_net,
    weight_bus_input_1 => delay_1_q_net,
    valid_bus_input_1 => enable_passthrough_case_1_y_net,
    hard_reset => switch_to_zero_y_net,
    pixel_bus_input_offset_0_2 => delay_108_q_net,
    pixel_bus_input_offset_0_3 => delay_114_q_net,
    pixel_bus_input_offset_0_4 => delay_116_q_net,
    pixel_bus_input_offset_0_5 => delay_118_q_net,
    pixel_bus_input_offset_0_6 => delay_98_q_net,
    pixel_bus_input_offset_0_7 => delay_100_q_net,
    pixel_bus_input_offset_0_8 => delay_102_q_net,
    pixel_bus_input_offset_0_9 => delay_111_q_net,
    pixel_bus_input_offset_0_10 => delay_104_q_net,
    pixel_bus_input_offset_0_11 => delay_106_q_net,
    pixel_bus_input_offset_0_12 => delay_109_q_net,
    pixel_bus_input_offset_1_2 => delay_2_q_net,
    pixel_bus_input_offset_1_3 => delay_4_q_net,
    pixel_bus_input_offset_1_4 => delay_6_q_net,
    pixel_bus_input_offset_1_5 => delay_8_q_net,
    pixel_bus_input_offset_1_6 => delay_10_q_net,
    pixel_bus_input_offset_1_7 => delay_12_q_net,
    pixel_bus_input_offset_1_8 => delay_14_q_net,
    pixel_bus_input_offset_1_9 => delay_23_q_net,
    pixel_bus_input_offset_1_10 => delay_16_q_net,
    pixel_bus_input_offset_1_11 => delay_18_q_net,
    pixel_bus_input_offset_1_12 => delay_20_q_net,
    pixel_bus_input_offset_2_2 => delay_36_q_net,
    pixel_bus_input_offset_2_3 => delay_42_q_net,
    pixel_bus_input_offset_2_4 => delay_44_q_net,
    pixel_bus_input_offset_2_5 => delay_46_q_net,
    pixel_bus_input_offset_2_6 => delay_26_q_net,
    pixel_bus_input_offset_2_7 => delay_28_q_net,
    pixel_bus_input_offset_2_8 => delay_30_q_net,
    pixel_bus_input_offset_2_9 => delay_39_q_net,
    pixel_bus_input_offset_2_10 => delay_32_q_net,
    pixel_bus_input_offset_2_11 => delay_34_q_net,
    pixel_bus_input_offset_2_12 => delay_37_q_net,
    pixel_bus_input_offset_3_2 => delay_60_q_net,
    pixel_bus_input_offset_3_3 => delay_66_q_net,
    pixel_bus_input_offset_3_4 => delay_68_q_net,
    pixel_bus_input_offset_3_5 => delay_70_q_net,
    pixel_bus_input_offset_3_6 => delay_50_q_net,
    pixel_bus_input_offset_3_7 => delay_52_q_net,
    pixel_bus_input_offset_3_8 => delay_54_q_net,
    pixel_bus_input_offset_3_9 => delay_63_q_net,
    pixel_bus_input_offset_3_10 => delay_56_q_net,
    pixel_bus_input_offset_3_11 => delay_58_q_net,
    pixel_bus_input_offset_3_12 => delay_61_q_net,
    pixel_bus_input_offset_4_2 => delay_84_q_net,
    pixel_bus_input_offset_4_3 => delay_90_q_net,
    pixel_bus_input_offset_4_4 => delay_92_q_net,
    pixel_bus_input_offset_4_5 => delay_94_q_net,
    pixel_bus_input_offset_4_6 => delay_74_q_net,
    pixel_bus_input_offset_4_7 => delay_76_q_net,
    pixel_bus_input_offset_4_8 => delay_78_q_net,
    pixel_bus_input_offset_4_9 => delay_87_q_net,
    pixel_bus_input_offset_4_10 => delay_80_q_net,
    pixel_bus_input_offset_4_11 => delay_82_q_net,
    pixel_bus_input_offset_4_12 => delay_85_q_net,
    weight_bus_input_2 => delay_3_q_net,
    weight_bus_input_3 => delay_5_q_net,
    weight_bus_input_4 => delay_7_q_net,
    weight_bus_input_5 => delay_9_q_net,
    weight_bus_input_6 => delay_11_q_net,
    weight_bus_input_7 => delay_13_q_net,
    weight_bus_input_8 => delay_15_q_net,
    weight_bus_input_9 => delay_24_q_net,
    weight_bus_input_10 => delay_17_q_net,
    weight_bus_input_11 => delay_19_q_net,
    weight_bus_input_12 => delay_21_q_net,
    weight_bus_input_13 => delay_25_q_net,
    weight_bus_input_14 => delay_41_q_net,
    weight_bus_input_15 => delay_43_q_net,
    weight_bus_input_16 => delay_45_q_net,
    weight_bus_input_17 => delay_47_q_net,
    weight_bus_input_18 => delay_27_q_net,
    weight_bus_input_19 => delay_29_q_net,
    weight_bus_input_20 => delay_31_q_net,
    weight_bus_input_21 => delay_40_q_net,
    weight_bus_input_22 => delay_33_q_net,
    weight_bus_input_23 => delay_35_q_net,
    weight_bus_input_24 => delay_38_q_net,
    weight_bus_input_25 => delay_49_q_net,
    weight_bus_input_26 => delay_65_q_net,
    weight_bus_input_27 => delay_67_q_net,
    weight_bus_input_28 => delay_69_q_net,
    weight_bus_input_29 => delay_71_q_net,
    weight_bus_input_30 => delay_51_q_net,
    weight_bus_input_31 => delay_53_q_net,
    weight_bus_input_32 => delay_55_q_net,
    weight_bus_input_33 => delay_64_q_net,
    weight_bus_input_34 => delay_57_q_net,
    weight_bus_input_35 => delay_59_q_net,
    weight_bus_input_36 => delay_62_q_net,
    weight_bus_input_37 => delay_73_q_net,
    weight_bus_input_38 => delay_89_q_net,
    weight_bus_input_39 => delay_91_q_net,
    weight_bus_input_40 => delay_93_q_net,
    weight_bus_input_41 => delay_95_q_net,
    weight_bus_input_42 => delay_75_q_net,
    weight_bus_input_43 => delay_77_q_net,
    weight_bus_input_44 => delay_79_q_net,
    weight_bus_input_45 => delay_88_q_net,
    weight_bus_input_46 => delay_81_q_net,
    weight_bus_input_47 => delay_83_q_net,
    weight_bus_input_48 => delay_86_q_net,
    weight_bus_input_49 => delay_97_q_net,
    weight_bus_input_50 => delay_113_q_net,
    weight_bus_input_51 => delay_115_q_net,
    weight_bus_input_52 => delay_117_q_net,
    weight_bus_input_53 => delay_119_q_net,
    weight_bus_input_54 => delay_99_q_net,
    weight_bus_input_55 => delay_101_q_net,
    weight_bus_input_56 => delay_103_q_net,
    weight_bus_input_57 => delay_112_q_net,
    weight_bus_input_58 => delay_105_q_net,
    weight_bus_input_59 => delay_107_q_net,
    weight_bus_input_60 => delay_110_q_net,
    weight_bus_input_61 => last_out_q_net,
    valid_bus_input_2 => enable_passthrough_case_0_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => accumulator_kernel_result_0_q_net_x7,
    valid_kernel_output => delay_enable_4_q_net_x6
  );
  subsystem : entity xil_defaultlib.mh_subsystem 
  port map (
    kernel_result_0 => accumulator_kernel_result_0_q_net_x6,
    kernel_result_valid_0 => delay_enable_4_q_net_x5,
    kernel_result_1 => accumulator_kernel_result_0_q_net_x5,
    kernel_result_valid_1 => delay_enable_4_q_net_x4,
    kernel_result_2 => accumulator_kernel_result_0_q_net_x4,
    kernel_result_valid_2 => delay_enable_4_q_net_x3,
    kernel_result_3 => accumulator_kernel_result_0_q_net_x3,
    kernel_result_valid_3 => delay_enable_4_q_net_x2,
    kernel_result_4 => accumulator_kernel_result_0_q_net_x2,
    kernel_result_valid_4 => delay_enable_4_q_net_x1,
    kernel_result_5 => accumulator_kernel_result_0_q_net_x1,
    kernel_result_valid_5 => delay_enable_4_q_net_x0,
    kernel_result_6 => accumulator_kernel_result_0_q_net_x0,
    kernel_result_valid_6 => delay_enable_4_q_net,
    kernel_result_7 => accumulator_kernel_result_0_q_net,
    kernel_result_valid_7 => delay_enable_4_q_net_x8,
    kernel_result_8 => accumulator_kernel_result_0_q_net_x8,
    kernel_result_valid_8 => delay_enable_4_q_net_x7,
    kernel_result_9 => accumulator_kernel_result_0_q_net_x7,
    kernel_result_valid_9 => delay_enable_4_q_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_result_output => output_or_block_y_net,
    kernel_result_output_valid => output_enable_y_net,
    kernel_result_array_position => kernel_result_array_offset_op_net,
    kernel_result_row_depth_position => kernel_result_array_offset1_op_net,
    finished_cube => switch_to_zero_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Frame Memory Controller
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_frame_memory_controller is
  port (
    x12_bit_data_in : in std_logic_vector( 12-1 downto 0 );
    enable_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_out_72_bits : out std_logic_vector( 72-1 downto 0 );
    data_out_ready : out std_logic_vector( 1-1 downto 0 );
    data_address_out : out std_logic_vector( 17-1 downto 0 );
    ram_bloack_sel_out : out std_logic_vector( 3-1 downto 0 );
    memory_is_full : out std_logic_vector( 1-1 downto 0 );
    new_frame_finished : out std_logic_vector( 1-1 downto 0 )
  );
end mh_frame_memory_controller;
architecture structural of mh_frame_memory_controller is 
  signal section_op_net : std_logic_vector( 8-1 downto 0 );
  signal or_offset_4_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal memory_full_delay_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal or_offset_5_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal zero_value1_y_net : std_logic_vector( 9-1 downto 0 );
  signal offset_fifo_0_full_net : std_logic;
  signal offset_fifo_3_full_net : std_logic;
  signal offset_fifo_1_full_net : std_logic;
  signal offset_fifo_4_full_net : std_logic;
  signal offset_fifo_2_full_net : std_logic;
  signal offset_fifo_5_full_net : std_logic;
  signal final_add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal add_ram_sel_delay_1_q_net : std_logic_vector( 3-1 downto 0 );
  signal clk_net : std_logic;
  signal memory_full_delay_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal and_input_delay_q_net : std_logic_vector( 12-1 downto 0 );
  signal and_input_delay2_q_net : std_logic_vector( 12-1 downto 0 );
  signal multiple_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_frame_and_section_s_net : std_logic_vector( 18-1 downto 0 );
  signal multiple_frame_p_net : std_logic_vector( 10-1 downto 0 );
  signal multiple_section_p_net : std_logic_vector( 17-1 downto 0 );
  signal mux_input_delay_q_net : std_logic_vector( 12-1 downto 0 );
  signal data_input_12_bit_net : std_logic_vector( 12-1 downto 0 );
  signal final_add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal add_offset_with_line_count_s_net : std_logic_vector( 17-1 downto 0 );
  signal ce_net : std_logic;
  signal multiple_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal write_enable_12_bit_net : std_logic_vector( 1-1 downto 0 );
  signal memory_full_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal and_ram_sel_delay_q_net : std_logic_vector( 3-1 downto 0 );
  signal check_for_new_line_op_net : std_logic_vector( 1-1 downto 0 );
  signal and_for_new_line_1099_check_y_net : std_logic_vector( 1-1 downto 0 );
  signal ram_block_determination_op_net : std_logic_vector( 3-1 downto 0 );
  signal check_for_new_frame_last_row_op_net : std_logic_vector( 1-1 downto 0 );
  signal add_ram_sel_delay_0_q_net : std_logic_vector( 3-1 downto 0 );
  signal add_line_delay_0_q_net : std_logic_vector( 7-1 downto 0 );
  signal multiple_ram_sel_delay_q_net : std_logic_vector( 3-1 downto 0 );
  signal check_new_frame_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_new_frame_last_pixel_op_net : std_logic_vector( 1-1 downto 0 );
  signal add_line_delay_1_q_net : std_logic_vector( 7-1 downto 0 );
  signal data_points_per_line_op_net : std_logic_vector( 7-1 downto 0 );
  signal and_for_new_line_y_net : std_logic_vector( 1-1 downto 0 );
  signal check_new_line_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_3_empty_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_1_empty_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal line_counter_op_net : std_logic_vector( 11-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 11-1 downto 0 );
  signal offset_fifo_4_empty_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 7-1 downto 0 );
  signal check_for_new_section_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_2_empty_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_0_empty_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_5_empty_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_last_pixel_on_ram_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_all_not_empty_y_net : std_logic_vector( 1-1 downto 0 );
  signal check_if_full_y_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_0_dout_net : std_logic_vector( 12-1 downto 0 );
  signal is_last_frame_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_3_dout_net : std_logic_vector( 12-1 downto 0 );
  signal offset_fifo_1_dout_net : std_logic_vector( 12-1 downto 0 );
  signal offset_fifo_5_dout_net : std_logic_vector( 12-1 downto 0 );
  signal check_if_full1_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_4_dout_net : std_logic_vector( 12-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 7-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 9-1 downto 0 );
  signal offset_fifo_2_dout_net : std_logic_vector( 12-1 downto 0 );
  signal concat_72_bit_packed_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal hold_up_read_out_op_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_5_op_net : std_logic_vector( 9-1 downto 0 );
  signal counter_compare_3_op_net : std_logic_vector( 9-1 downto 0 );
  signal enable_offset_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_offset_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_4_op_net : std_logic_vector( 9-1 downto 0 );
  signal enable_offset_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_1_op_net : std_logic_vector( 9-1 downto 0 );
  signal counter_compare_2_op_net : std_logic_vector( 9-1 downto 0 );
  signal counter_compare_0_op_net : std_logic_vector( 9-1 downto 0 );
  signal convert_to_bool_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_2_cycle_enable_to_1_cycle_op_net : std_logic_vector( 2-1 downto 0 );
  signal enable_offset_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_offset_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal offset_2_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_3_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal data_points_op_net : std_logic_vector( 9-1 downto 0 );
  signal mux_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_0_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_4_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_5_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_1_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal enable_offset_5_y_net : std_logic_vector( 1-1 downto 0 );
  signal frame_op_net : std_logic_vector( 3-1 downto 0 );
  signal mux_delay_we_fifo_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal last_value_to_pack_op_net : std_logic_vector( 9-1 downto 0 );
  signal impossible_value_op_net : std_logic_vector( 9-1 downto 0 );
  signal mux_delay_input_q_net : std_logic_vector( 12-1 downto 0 );
  signal mux_enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_4_check1_op_net : std_logic_vector( 1-1 downto 0 );
  signal zero_out_op_net : std_logic_vector( 12-1 downto 0 );
  signal mux_delay_we_fifo_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_delay_we_fifo_3_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_zero_value_or_input_data_y_net : std_logic_vector( 12-1 downto 0 );
  signal mux_delay_we_fifo_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mass_enable_offset_y_net : std_logic_vector( 1-1 downto 0 );
begin
  data_out_72_bits <= final_add_data_out_delay_q_net;
  data_out_ready <= final_add_enable_delay_q_net;
  data_address_out <= add_offset_with_line_count_s_net;
  ram_bloack_sel_out <= add_ram_sel_delay_1_q_net;
  memory_is_full <= memory_full_delay_1_q_net;
  new_frame_finished <= memory_full_delay_2_q_net;
  data_input_12_bit_net <= x12_bit_data_in;
  write_enable_12_bit_net <= enable_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  and_input_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_input_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => and_input_delay_q_net
  );
  and_input_delay2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => and_input_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => and_input_delay2_q_net
  );
  add_data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => multiple_data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_data_out_delay_q_net
  );
  add_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => multiple_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_enable_delay_q_net
  );
  add_frame_and_section : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 10,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 17,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "mh_c_addsub_v12_0_i7",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 18,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => multiple_frame_p_net,
    b => multiple_section_p_net,
    clk => clk_net,
    ce => ce_net,
    s => add_frame_and_section_s_net
  );
  add_line_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 7
  )
  port map (
    en => '1',
    rst => '0',
    d => data_points_per_line_op_net,
    clk => clk_net,
    ce => ce_net,
    q => add_line_delay_0_q_net
  );
  add_line_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 7
  )
  port map (
    en => '1',
    rst => '0',
    d => add_line_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_line_delay_1_q_net
  );
  add_offset_with_line_count : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 7,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "mh_c_addsub_v12_0_i8",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => add_line_delay_1_q_net,
    b => add_frame_and_section_s_net,
    clk => clk_net,
    ce => ce_net,
    s => add_offset_with_line_count_s_net
  );
  add_ram_sel_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => multiple_ram_sel_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_ram_sel_delay_0_q_net
  );
  add_ram_sel_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => add_ram_sel_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_ram_sel_delay_1_q_net
  );
  and_ram_sel_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => ram_block_determination_op_net,
    clk => clk_net,
    ce => ce_net,
    q => and_ram_sel_delay_q_net
  );
  and_for_new_line : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => check_for_new_line_op_net,
    d1 => check_new_line_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => and_for_new_line_y_net
  );
  and_for_new_line_1099_check : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => check_for_new_frame_last_row_op_net,
    d1 => check_new_frame_enable_delay_q_net,
    d2 => check_for_new_frame_last_pixel_op_net,
    clk => clk_net,
    ce => ce_net,
    y => and_for_new_line_1099_check_y_net
  );
  check_for_all_not_empty : entity xil_defaultlib.sysgen_logical_8143a363af 
  port map (
    clr => '0',
    d0 => offset_fifo_5_empty_net,
    d1 => offset_fifo_4_empty_net,
    d2 => offset_fifo_3_empty_net,
    d3 => offset_fifo_2_empty_net,
    d4 => offset_fifo_1_empty_net,
    d5 => offset_fifo_0_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => check_for_all_not_empty_y_net
  );
  check_for_new_frame_last_pixel : entity xil_defaultlib.sysgen_relational_66ac941b9b 
  port map (
    clr => '0',
    a => data_points_per_line_op_net,
    b => constant2_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => check_for_new_frame_last_pixel_op_net
  );
  check_new_frame_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    q => check_new_frame_enable_delay_q_net
  );
  check_new_line_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    q => check_new_line_delay_q_net
  );
  check_for_new_frame_last_row : entity xil_defaultlib.sysgen_relational_22128290a8 
  port map (
    clr => '0',
    a => line_counter_op_net,
    b => constant4_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => check_for_new_frame_last_row_op_net
  );
  check_for_last_pixel_on_ram_4 : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => check_for_new_section_op_net,
    d1 => check_new_frame_enable_delay_q_net,
    d2 => check_for_new_frame_last_pixel_op_net,
    clk => clk_net,
    ce => ce_net,
    y => check_for_last_pixel_on_ram_4_y_net
  );
  check_for_new_line : entity xil_defaultlib.sysgen_relational_66ac941b9b 
  port map (
    clr => '0',
    a => data_points_per_line_op_net,
    b => constant2_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => check_for_new_line_op_net
  );
  check_for_new_section : entity xil_defaultlib.sysgen_relational_4b66a02210 
  port map (
    clr => '0',
    a => constant6_op_net,
    b => ram_block_determination_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => check_for_new_section_op_net
  );
  check_if_full : entity xil_defaultlib.sysgen_logical_f8bf58b41a 
  port map (
    clr => '0',
    d0 => check_for_new_frame_last_row_op_net,
    d1 => check_for_new_frame_last_pixel_op_net,
    d2 => check_new_frame_enable_delay_q_net,
    d3 => is_last_frame_op_net,
    clk => clk_net,
    ce => ce_net,
    y => check_if_full_y_net
  );
  check_if_full1 : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => check_for_new_frame_last_row_op_net,
    d1 => check_for_new_frame_last_pixel_op_net,
    d2 => check_new_frame_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => check_if_full1_y_net
  );
  concat_72_bit_packed_value : entity xil_defaultlib.sysgen_concat_e690ad1743 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => offset_fifo_5_dout_net,
    in1 => offset_fifo_4_dout_net,
    in2 => offset_fifo_3_dout_net,
    in3 => offset_fifo_2_dout_net,
    in4 => offset_fifo_1_dout_net,
    in5 => offset_fifo_0_dout_net,
    y => concat_72_bit_packed_value_y_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_6b755964f8 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_e7009a7f9c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_30acb293d3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_44db6fe362 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  convert_2_cycle_enable_to_1_cycle : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    rst => "0",
    clr => '0',
    en => check_for_all_not_empty_y_net,
    clk => clk_net,
    ce => ce_net,
    op => convert_2_cycle_enable_to_1_cycle_op_net
  );
  convert_to_bool : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 3,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => hold_up_read_out_op_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_to_bool_dout_net
  );
  convert_to_bool_x0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 2,
    y_width => 1
  )
  port map (
    x => convert_2_cycle_enable_to_1_cycle_op_net,
    y => convert_to_bool_y_net
  );
  counter_compare_0 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 396,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i4",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_offset_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_0_op_net
  );
  counter_compare_1 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 397,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i5",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_offset_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_1_op_net
  );
  counter_compare_2 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 398,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i6",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_offset_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_2_op_net
  );
  counter_compare_3 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 399,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i7",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_offset_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_3_op_net
  );
  counter_compare_4 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 394,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i8",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_offset_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_4_op_net
  );
  counter_compare_5 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 395,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i9",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_offset_5_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_5_op_net
  );
  data_points : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 399,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i10",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => write_enable_12_bit_net,
    clk => clk_net,
    ce => ce_net,
    op => data_points_op_net
  );
  data_points_per_line : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 66,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i0",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    rst => "0",
    clr => '0',
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => data_points_per_line_op_net
  );
  enable_offset_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_0_check_op_net,
    d1 => mux_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_offset_0_y_net
  );
  enable_offset_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_1_check_op_net,
    d1 => mux_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_offset_1_y_net
  );
  enable_offset_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_2_check_op_net,
    d1 => mux_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_offset_2_y_net
  );
  enable_offset_3 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_3_check_op_net,
    d1 => mux_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_offset_3_y_net
  );
  enable_offset_4 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_4_check_op_net,
    d1 => mux_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_offset_4_y_net
  );
  enable_offset_5 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_5_check_op_net,
    d1 => mux_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_offset_5_y_net
  );
  fifo_delay_enable : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_to_bool_y_net,
    clk => clk_net,
    ce => ce_net,
    q => fifo_delay_enable_q_net
  );
  final_add_data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => add_data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => final_add_data_out_delay_q_net
  );
  final_add_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => add_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => final_add_enable_delay_q_net
  );
  frame : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 4,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i11",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 3
  )
  port map (
    rst => "0",
    clr => '0',
    en => and_for_new_line_1099_check_y_net,
    clk => clk_net,
    ce => ce_net,
    op => frame_op_net
  );
  hold_up_read_out : entity xil_defaultlib.sysgen_counter_27d1542d0d 
  port map (
    clr => '0',
    load => check_if_full_y_net,
    din => constant7_op_net,
    en => check_if_full_y_net,
    clk => clk_net,
    ce => ce_net,
    op => hold_up_read_out_op_net
  );
  impossible_value : entity xil_defaultlib.sysgen_constant_a034db8e06 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => impossible_value_op_net
  );
  is_last_frame : entity xil_defaultlib.sysgen_relational_4b66a02210 
  port map (
    clr => '0',
    a => frame_op_net,
    b => constant6_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => is_last_frame_op_net
  );
  last_value_to_pack : entity xil_defaultlib.sysgen_constant_40850aac15 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => last_value_to_pack_op_net
  );
  line_counter : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 1099,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i12",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 11
  )
  port map (
    rst => "0",
    clr => '0',
    en => and_for_new_line_y_net,
    clk => clk_net,
    ce => ce_net,
    op => line_counter_op_net
  );
  mux_delay_input : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => and_input_delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_delay_input_q_net
  );
  mux_delay_we_fifo_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_offset_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_delay_we_fifo_0_q_net
  );
  mux_delay_we_fifo_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_offset_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_delay_we_fifo_1_q_net
  );
  mux_delay_we_fifo_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_offset_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_delay_we_fifo_2_q_net
  );
  mux_delay_we_fifo_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => enable_offset_3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_delay_we_fifo_3_q_net
  );
  mux_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay_q_net
  );
  mux_enable_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => write_enable_12_bit_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_enable_delay1_q_net
  );
  mux_input_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => data_input_12_bit_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_input_delay_q_net
  );
  mux_zero_value_or_input_data : entity xil_defaultlib.sysgen_mux_98805571d1 
  port map (
    clr => '0',
    sel => mass_enable_offset_y_net,
    d0 => and_input_delay2_q_net,
    d1 => zero_out_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_zero_value_or_input_data_y_net
  );
  mass_enable_offset : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => offset_4_check1_op_net,
    d1 => mux_enable_delay_q_net,
    d2 => offset_3_check_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mass_enable_offset_y_net
  );
  memory_full_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_to_bool_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => memory_full_delay_0_q_net
  );
  memory_full_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => memory_full_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => memory_full_delay_1_q_net
  );
  memory_full_delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 6,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => check_if_full1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => memory_full_delay_2_q_net
  );
  multiple_data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => concat_72_bit_packed_value_y_net,
    clk => clk_net,
    ce => ce_net,
    q => multiple_data_out_delay_q_net
  );
  multiple_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    q => multiple_enable_delay_q_net
  );
  multiple_frame : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 7,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 3,
    c_a_type => 1,
    c_a_width => 7,
    c_b_type => 1,
    c_b_width => 3,
    c_baat => 7,
    c_output_width => 10,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i1",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 10,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => constant3_op_net,
    b => frame_op_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => multiple_frame_p_net
  );
  multiple_ram_sel_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => and_ram_sel_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => multiple_ram_sel_delay_q_net
  );
  multiple_section : entity xil_defaultlib.mh_xlmult 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 9,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 8,
    c_a_type => 1,
    c_a_width => 9,
    c_b_type => 1,
    c_b_width => 8,
    c_baat => 9,
    c_output_width => 17,
    c_type => 1,
    core_name0 => "mh_mult_gen_v12_0_i2",
    extra_registers => 0,
    multsign => 1,
    overflow => 1,
    p_arith => xlUnsigned,
    p_bin_pt => 0,
    p_width => 17,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => constant5_op_net,
    b => section_op_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => multiple_section_p_net
  );
  or_offset_4_enable : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => mass_enable_offset_y_net,
    d1 => enable_offset_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => or_offset_4_enable_y_net
  );
  or_offset_5_enable : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => enable_offset_5_y_net,
    d1 => mass_enable_offset_y_net,
    clk => clk_net,
    ce => ce_net,
    y => or_offset_5_enable_y_net
  );
  offset_0_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => zero_value1_y_net,
    b => counter_compare_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_0_check_op_net
  );
  offset_1_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => zero_value1_y_net,
    b => counter_compare_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_1_check_op_net
  );
  offset_2_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => zero_value1_y_net,
    b => counter_compare_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_2_check_op_net
  );
  offset_3_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => zero_value1_y_net,
    b => counter_compare_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_3_check_op_net
  );
  offset_4_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => zero_value1_y_net,
    b => counter_compare_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_4_check_op_net
  );
  offset_4_check1 : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => last_value_to_pack_op_net,
    b => zero_value1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_4_check1_op_net
  );
  offset_5_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => zero_value1_y_net,
    b => counter_compare_5_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_5_check_op_net
  );
  offset_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i1",
    data_count_width => 4,
    data_width => 12,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => mux_delay_input_q_net,
    we => mux_delay_we_fifo_0_q_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_0_dout_net,
    empty => offset_fifo_0_empty_net(0),
    full => offset_fifo_0_full_net
  );
  offset_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i1",
    data_count_width => 4,
    data_width => 12,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => mux_delay_input_q_net,
    we => mux_delay_we_fifo_1_q_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_1_dout_net,
    empty => offset_fifo_1_empty_net(0),
    full => offset_fifo_1_full_net
  );
  offset_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i1",
    data_count_width => 4,
    data_width => 12,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => mux_delay_input_q_net,
    we => mux_delay_we_fifo_2_q_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_2_dout_net,
    empty => offset_fifo_2_empty_net(0),
    full => offset_fifo_2_full_net
  );
  offset_fifo_3 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i1",
    data_count_width => 4,
    data_width => 12,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => mux_delay_input_q_net,
    we => mux_delay_we_fifo_3_q_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_3_dout_net,
    empty => offset_fifo_3_empty_net(0),
    full => offset_fifo_3_full_net
  );
  offset_fifo_4 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i1",
    data_count_width => 4,
    data_width => 12,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => mux_zero_value_or_input_data_y_net,
    we => or_offset_4_enable_y_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_4_dout_net,
    empty => offset_fifo_4_empty_net(0),
    full => offset_fifo_4_full_net
  );
  offset_fifo_5 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i1",
    data_count_width => 4,
    data_width => 12,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => mux_zero_value_or_input_data_y_net,
    we => or_offset_5_enable_y_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_5_dout_net,
    empty => offset_fifo_5_empty_net(0),
    full => offset_fifo_5_full_net
  );
  ram_block_determination : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 4,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i11",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 3
  )
  port map (
    rst => "0",
    clr => '0',
    en => and_for_new_line_y_net,
    clk => clk_net,
    ce => ce_net,
    op => ram_block_determination_op_net
  );
  section : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 219,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i13",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    rst => "0",
    clr => '0',
    en => check_for_last_pixel_on_ram_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => section_op_net
  );
  zero_out : entity xil_defaultlib.sysgen_constant_bdf9cca84c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => zero_out_op_net
  );
  zero_value1 : entity xil_defaultlib.sysgen_mux_044d346e3b 
  port map (
    clr => '0',
    sel => write_enable_12_bit_net,
    d0 => impossible_value_op_net,
    d1 => data_points_op_net,
    clk => clk_net,
    ce => ce_net,
    y => zero_value1_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Kernel Memory Controller
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_memory_controller is
  port (
    x18_bit_data_in : in std_logic_vector( 18-1 downto 0 );
    enable_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_out_72_bits : out std_logic_vector( 72-1 downto 0 );
    data_out_ready : out std_logic_vector( 1-1 downto 0 );
    data_address_out : out std_logic_vector( 9-1 downto 0 );
    ram_block_sel_out : out std_logic_vector( 3-1 downto 0 );
    memory_is_full : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_memory_controller;
architecture structural of mh_kernel_memory_controller is 
  signal ce_net : std_logic;
  signal multiple_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal final_add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal add_ram_sel_delay_1_q_net : std_logic_vector( 3-1 downto 0 );
  signal final_add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal multiple_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_18_bit_net : std_logic_vector( 18-1 downto 0 );
  signal data_points_per_line_op_net : std_logic_vector( 9-1 downto 0 );
  signal memory_full_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal data_out_delay_q_net : std_logic_vector( 9-1 downto 0 );
  signal add_line_delay_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal data_enable_18_bit_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_0_empty_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_3_empty_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_new_section_op_net : std_logic_vector( 1-1 downto 0 );
  signal check_new_line_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_2_empty_net : std_logic_vector( 1-1 downto 0 );
  signal add_line_delay_1_q_net : std_logic_vector( 9-1 downto 0 );
  signal check_for_all_not_empty_y_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_1_empty_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_new_line_op_net : std_logic_vector( 1-1 downto 0 );
  signal add_ram_sel_delay_0_q_net : std_logic_vector( 3-1 downto 0 );
  signal and_for_new_section_y_net : std_logic_vector( 1-1 downto 0 );
  signal multiple_ram_sel_delay_q_net : std_logic_vector( 3-1 downto 0 );
  signal check_new_for_ands_q_net : std_logic_vector( 1-1 downto 0 );
  signal and_for_new_line_y_net : std_logic_vector( 1-1 downto 0 );
  signal compare_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 3-1 downto 0 );
  signal offset_fifo_0_dout_net : std_logic_vector( 18-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 1-1 downto 0 );
  signal check_if_full_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat_72_bit_packed_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal mux_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 12-1 downto 0 );
  signal offset_fifo_3_dout_net : std_logic_vector( 18-1 downto 0 );
  signal offset_fifo_2_dout_net : std_logic_vector( 18-1 downto 0 );
  signal offset_fifo_1_dout_net : std_logic_vector( 18-1 downto 0 );
  signal ram_block_determination_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 9-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_2_op_net : std_logic_vector( 9-1 downto 0 );
  signal data_points_op_net : std_logic_vector( 9-1 downto 0 );
  signal write_enable_offset_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_1_op_net : std_logic_vector( 9-1 downto 0 );
  signal convert_2_cycle_enable_to_1_cycle_op_net : std_logic_vector( 2-1 downto 0 );
  signal hold_up_read_out_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_enable_offset_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_enable_offset_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_3_op_net : std_logic_vector( 9-1 downto 0 );
  signal counter_compare_0_op_net : std_logic_vector( 9-1 downto 0 );
  signal write_enable_offset_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_write_enable_and_q_net : std_logic_vector( 18-1 downto 0 );
  signal memory_full_delay_0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_write_enable_checking_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_write_enable_mux_q_net : std_logic_vector( 18-1 downto 0 );
  signal offset_1_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_0_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_2_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal offset_3_check_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 9-1 downto 0 );
  signal offset_fifo_0_full_net : std_logic;
  signal offset_fifo_2_full_net : std_logic;
  signal offset_fifo_3_full_net : std_logic;
  signal offset_fifo_1_full_net : std_logic;
begin
  data_out_72_bits <= final_add_data_out_delay_q_net;
  data_out_ready <= final_add_enable_delay_q_net;
  data_address_out <= data_out_delay_q_net;
  ram_block_sel_out <= add_ram_sel_delay_1_q_net;
  memory_is_full <= memory_full_delay_1_q_net;
  data_in_18_bit_net <= x18_bit_data_in;
  data_enable_18_bit_net <= enable_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  add_data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => multiple_data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_data_out_delay_q_net
  );
  add_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => multiple_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_enable_delay_q_net
  );
  add_line_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => data_points_per_line_op_net,
    clk => clk_net,
    ce => ce_net,
    q => add_line_delay_0_q_net
  );
  add_line_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => add_line_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_line_delay_1_q_net
  );
  add_ram_sel_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => multiple_ram_sel_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_ram_sel_delay_0_q_net
  );
  add_ram_sel_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => add_ram_sel_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => add_ram_sel_delay_1_q_net
  );
  and_for_new_line : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => check_for_new_line_op_net,
    d1 => check_new_line_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => and_for_new_line_y_net
  );
  and_for_new_section : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => check_new_line_delay_q_net,
    d1 => check_for_new_section_op_net,
    clk => clk_net,
    ce => ce_net,
    y => and_for_new_section_y_net
  );
  check_for_all_not_empty : entity xil_defaultlib.sysgen_logical_e1ed02b118 
  port map (
    clr => '0',
    d0 => offset_fifo_2_empty_net,
    d1 => offset_fifo_3_empty_net,
    d2 => offset_fifo_1_empty_net,
    d3 => offset_fifo_0_empty_net,
    clk => clk_net,
    ce => ce_net,
    y => check_for_all_not_empty_y_net
  );
  check_new_for_ands : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => check_new_line_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => check_new_for_ands_q_net
  );
  check_new_line_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    q => check_new_line_delay_q_net
  );
  check_for_new_line : entity xil_defaultlib.sysgen_relational_543814c385 
  port map (
    clr => '0',
    a => data_points_per_line_op_net,
    b => constant2_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => check_for_new_line_op_net
  );
  check_for_new_section : entity xil_defaultlib.sysgen_relational_4b66a02210 
  port map (
    clr => '0',
    a => ram_block_determination_op_net,
    b => constant6_op_net,
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => check_for_new_section_op_net
  );
  check_if_full : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => and_for_new_line_y_net,
    d1 => check_new_for_ands_q_net,
    d2 => and_for_new_section_y_net,
    clk => clk_net,
    ce => ce_net,
    y => check_if_full_y_net
  );
  compare_delay_enable : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => mux_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_delay_enable_q_net
  );
  concat_72_bit_packed_value : entity xil_defaultlib.sysgen_concat_dcc3502f5b 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => offset_fifo_3_dout_net,
    in1 => offset_fifo_2_dout_net,
    in2 => offset_fifo_1_dout_net,
    in3 => offset_fifo_0_dout_net,
    y => concat_72_bit_packed_value_y_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_a034db8e06 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_2a0c3f2acd 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  convert_2_cycle_enable_to_1_cycle : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    rst => "0",
    clr => '0',
    en => check_for_all_not_empty_y_net,
    clk => clk_net,
    ce => ce_net,
    op => convert_2_cycle_enable_to_1_cycle_op_net
  );
  convert_to_bool : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 3,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => hold_up_read_out_op_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_to_bool_dout_net
  );
  convert_to_bool_x0 : entity xil_defaultlib.mh_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 2,
    y_width => 1
  )
  port map (
    x => convert_2_cycle_enable_to_1_cycle_op_net,
    y => convert_to_bool_y_net
  );
  counter_compare_0 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 396,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i14",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => write_enable_offset_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_0_op_net
  );
  counter_compare_1 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 397,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i15",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => write_enable_offset_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_1_op_net
  );
  counter_compare_2 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 398,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i16",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => write_enable_offset_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_2_op_net
  );
  counter_compare_3 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 399,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i17",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => write_enable_offset_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_compare_3_op_net
  );
  data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => add_line_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => data_out_delay_q_net
  );
  data_points : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 399,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i10",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => data_enable_18_bit_net,
    clk => clk_net,
    ce => ce_net,
    op => data_points_op_net
  );
  data_points_per_line : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 499,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i10",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    op => data_points_per_line_op_net
  );
  delay_write_enable_and : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_write_enable_checking_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_write_enable_and_q_net
  );
  delay_write_enable_checking : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_write_enable_mux_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_write_enable_checking_q_net
  );
  delay_write_enable_mux : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => data_in_18_bit_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_write_enable_mux_q_net
  );
  fifo_delay_enable : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_to_bool_y_net,
    clk => clk_net,
    ce => ce_net,
    q => fifo_delay_enable_q_net
  );
  final_add_data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => add_data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => final_add_data_out_delay_q_net
  );
  final_add_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => add_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => final_add_enable_delay_q_net
  );
  hold_up_read_out : entity xil_defaultlib.sysgen_counter_27d1542d0d 
  port map (
    clr => '0',
    load => check_if_full_y_net,
    din => constant7_op_net,
    en => check_if_full_y_net,
    clk => clk_net,
    ce => ce_net,
    op => hold_up_read_out_op_net
  );
  mux_delay_enable : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => data_enable_18_bit_net,
    clk => clk_net,
    ce => ce_net,
    q => mux_delay_enable_q_net
  );
  memory_full_delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_to_bool_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => memory_full_delay_0_q_net
  );
  memory_full_delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => memory_full_delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => memory_full_delay_1_q_net
  );
  multiple_data_out_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => concat_72_bit_packed_value_y_net,
    clk => clk_net,
    ce => ce_net,
    q => multiple_data_out_delay_q_net
  );
  multiple_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => fifo_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    q => multiple_enable_delay_q_net
  );
  multiple_ram_sel_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => ram_block_determination_op_net,
    clk => clk_net,
    ce => ce_net,
    q => multiple_ram_sel_delay_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_044d346e3b 
  port map (
    clr => '0',
    sel => data_enable_18_bit_net,
    d0 => constant1_op_net,
    d1 => data_points_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  offset_0_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => mux_y_net,
    b => counter_compare_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_0_check_op_net
  );
  offset_1_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => mux_y_net,
    b => counter_compare_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_1_check_op_net
  );
  offset_2_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => mux_y_net,
    b => counter_compare_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_2_check_op_net
  );
  offset_3_check : entity xil_defaultlib.sysgen_relational_7e53eec433 
  port map (
    clr => '0',
    a => mux_y_net,
    b => counter_compare_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => offset_3_check_op_net
  );
  offset_fifo_0 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i2",
    data_count_width => 4,
    data_width => 18,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => delay_write_enable_and_q_net,
    we => write_enable_offset_0_y_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_0_dout_net,
    empty => offset_fifo_0_empty_net(0),
    full => offset_fifo_0_full_net
  );
  offset_fifo_1 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i2",
    data_count_width => 4,
    data_width => 18,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => delay_write_enable_and_q_net,
    we => write_enable_offset_1_y_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_1_dout_net,
    empty => offset_fifo_1_empty_net(0),
    full => offset_fifo_1_full_net
  );
  offset_fifo_2 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i2",
    data_count_width => 4,
    data_width => 18,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => delay_write_enable_and_q_net,
    we => write_enable_offset_2_y_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_2_dout_net,
    empty => offset_fifo_2_empty_net(0),
    full => offset_fifo_2_full_net
  );
  offset_fifo_3 : entity xil_defaultlib.mh_xlfifogen_u 
  generic map (
    core_name0 => "mh_fifo_generator_i2",
    data_count_width => 4,
    data_width => 18,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 4
  )
  port map (
    en => '1',
    rst => '0',
    din => delay_write_enable_and_q_net,
    we => write_enable_offset_3_y_net(0),
    re => convert_to_bool_y_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => offset_fifo_3_dout_net,
    empty => offset_fifo_3_empty_net(0),
    full => offset_fifo_3_full_net
  );
  ram_block_determination : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 4,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i11",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 3
  )
  port map (
    rst => "0",
    clr => '0',
    en => and_for_new_line_y_net,
    clk => clk_net,
    ce => ce_net,
    op => ram_block_determination_op_net
  );
  write_enable_offset_0 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_0_check_op_net,
    d1 => compare_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_enable_offset_0_y_net
  );
  write_enable_offset_1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_1_check_op_net,
    d1 => compare_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_enable_offset_1_y_net
  );
  write_enable_offset_2 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_2_check_op_net,
    d1 => compare_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_enable_offset_2_y_net
  );
  write_enable_offset_3 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => offset_3_check_op_net,
    d1 => compare_delay_enable_q_net,
    clk => clk_net,
    ce => ce_net,
    y => write_enable_offset_3_y_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Kernel Memory Subsystem/RAM Selector 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_ram_selector_0 is
  port (
    data_in : in std_logic_vector( 9-1 downto 0 );
    ram_select : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_ram_0 : out std_logic_vector( 9-1 downto 0 );
    out_ram_1 : out std_logic_vector( 9-1 downto 0 );
    out_ram_2 : out std_logic_vector( 9-1 downto 0 );
    out_ram_3 : out std_logic_vector( 9-1 downto 0 );
    out_ram_4 : out std_logic_vector( 9-1 downto 0 )
  );
end mh_ram_selector_0;
architecture structural of mh_ram_selector_0 is 
  signal sel_ram_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 9-1 downto 0 );
  signal clk_net : std_logic;
  signal line_out_ram_1_y_net : std_logic_vector( 9-1 downto 0 );
  signal sel_ram_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_4_y_net : std_logic_vector( 9-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 9-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_q_net : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_1_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_3_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_4_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_0_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_2_op_net : std_logic_vector( 3-1 downto 0 );
begin
  out_ram_0 <= line_out_ram_0_y_net;
  out_ram_1 <= line_out_ram_1_y_net;
  out_ram_2 <= line_out_ram_2_y_net;
  out_ram_3 <= line_out_ram_3_y_net;
  out_ram_4 <= line_out_ram_4_y_net;
  delay_2_q_net <= data_in;
  delay_3_q_net <= ram_select;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  line_out_ram_0 : entity xil_defaultlib.sysgen_mux_2ddf659e9e 
  port map (
    clr => '0',
    sel => sel_ram_0_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_0_y_net
  );
  line_out_ram_1 : entity xil_defaultlib.sysgen_mux_2ddf659e9e 
  port map (
    clr => '0',
    sel => sel_ram_1_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_1_y_net
  );
  line_out_ram_2 : entity xil_defaultlib.sysgen_mux_2ddf659e9e 
  port map (
    clr => '0',
    sel => sel_ram_2_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_2_y_net
  );
  line_out_ram_3 : entity xil_defaultlib.sysgen_mux_2ddf659e9e 
  port map (
    clr => '0',
    sel => sel_ram_3_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_3_y_net
  );
  line_out_ram_4 : entity xil_defaultlib.sysgen_mux_2ddf659e9e 
  port map (
    clr => '0',
    sel => sel_ram_4_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_4_y_net
  );
  sel_ram_0 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_0_op_net
  );
  sel_ram_1 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_1_op_net
  );
  sel_ram_2 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_2_op_net
  );
  sel_ram_3 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_3_op_net
  );
  sel_ram_4 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_4_op_net
  );
  sel_value_ram_0 : entity xil_defaultlib.sysgen_constant_28e1aa0294 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_0_op_net
  );
  sel_value_ram_1 : entity xil_defaultlib.sysgen_constant_031f960172 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_1_op_net
  );
  sel_value_ram_2 : entity xil_defaultlib.sysgen_constant_15681d4665 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_2_op_net
  );
  sel_value_ram_3 : entity xil_defaultlib.sysgen_constant_c571582d8a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_3_op_net
  );
  sel_value_ram_4 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_4_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Kernel Memory Subsystem/RAM Selector 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_ram_selector_1 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    ram_select : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_ram_0 : out std_logic_vector( 72-1 downto 0 );
    out_ram_1 : out std_logic_vector( 72-1 downto 0 );
    out_ram_2 : out std_logic_vector( 72-1 downto 0 );
    out_ram_3 : out std_logic_vector( 72-1 downto 0 );
    out_ram_4 : out std_logic_vector( 72-1 downto 0 )
  );
end mh_ram_selector_1;
architecture structural of mh_ram_selector_1 is 
  signal clk_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 72-1 downto 0 );
  signal sel_ram_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_4_y_net : std_logic_vector( 72-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_1_y_net : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal sel_value_ram_3_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_2_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_1_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_0_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_4_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_4_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out_ram_0 <= line_out_ram_0_y_net;
  out_ram_1 <= line_out_ram_1_y_net;
  out_ram_2 <= line_out_ram_2_y_net;
  out_ram_3 <= line_out_ram_3_y_net;
  out_ram_4 <= line_out_ram_4_y_net;
  delay_0_q_net <= data_in;
  delay_3_q_net <= ram_select;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  line_out_ram_0 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_0_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_0_y_net
  );
  line_out_ram_1 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_1_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_1_y_net
  );
  line_out_ram_2 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_2_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_2_y_net
  );
  line_out_ram_3 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_3_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_3_y_net
  );
  line_out_ram_4 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_4_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_4_y_net
  );
  sel_ram_0 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_0_op_net
  );
  sel_ram_1 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_1_op_net
  );
  sel_ram_2 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_2_op_net
  );
  sel_ram_3 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_3_op_net
  );
  sel_ram_4 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_4_op_net
  );
  sel_value_ram_0 : entity xil_defaultlib.sysgen_constant_28e1aa0294 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_0_op_net
  );
  sel_value_ram_1 : entity xil_defaultlib.sysgen_constant_031f960172 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_1_op_net
  );
  sel_value_ram_2 : entity xil_defaultlib.sysgen_constant_15681d4665 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_2_op_net
  );
  sel_value_ram_3 : entity xil_defaultlib.sysgen_constant_c571582d8a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_3_op_net
  );
  sel_value_ram_4 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_4_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Kernel Memory Subsystem/RAM Selector 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_ram_selector_2_x0 is
  port (
    data_in : in std_logic_vector( 1-1 downto 0 );
    ram_select : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_ram_0 : out std_logic_vector( 1-1 downto 0 );
    out_ram_1 : out std_logic_vector( 1-1 downto 0 );
    out_ram_2 : out std_logic_vector( 1-1 downto 0 );
    out_ram_3 : out std_logic_vector( 1-1 downto 0 );
    out_ram_4 : out std_logic_vector( 1-1 downto 0 )
  );
end mh_ram_selector_2_x0;
architecture structural of mh_ram_selector_2_x0 is 
  signal sel_ram_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal line_out_ram_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_2_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_4_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_1_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_0_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_3_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_2_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out_ram_0 <= line_out_ram_0_y_net;
  out_ram_1 <= line_out_ram_1_y_net;
  out_ram_2 <= line_out_ram_2_y_net;
  out_ram_3 <= line_out_ram_3_y_net;
  out_ram_4 <= line_out_ram_4_y_net;
  delay_1_q_net <= data_in;
  delay_3_q_net <= ram_select;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  line_out_ram_0 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_0_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_0_y_net
  );
  line_out_ram_1 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_1_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_1_y_net
  );
  line_out_ram_2 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_2_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_2_y_net
  );
  line_out_ram_3 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_3_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_3_y_net
  );
  line_out_ram_4 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_4_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_4_y_net
  );
  sel_ram_0 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_0_op_net
  );
  sel_ram_1 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_1_op_net
  );
  sel_ram_2 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_2_op_net
  );
  sel_ram_3 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_3_op_net
  );
  sel_ram_4 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_4_op_net
  );
  sel_value_ram_0 : entity xil_defaultlib.sysgen_constant_28e1aa0294 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_0_op_net
  );
  sel_value_ram_1 : entity xil_defaultlib.sysgen_constant_031f960172 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_1_op_net
  );
  sel_value_ram_2 : entity xil_defaultlib.sysgen_constant_15681d4665 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_2_op_net
  );
  sel_value_ram_3 : entity xil_defaultlib.sysgen_constant_c571582d8a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_3_op_net
  );
  sel_value_ram_4 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_4_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Kernel Memory Subsystem
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_memory_subsystem is
  port (
    read_address : in std_logic_vector( 9-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    write_address : in std_logic_vector( 9-1 downto 0 );
    write_data_to_ram_sel : in std_logic_vector( 3-1 downto 0 );
    data_to_write : in std_logic_vector( 72-1 downto 0 );
    write_enable : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ram_0_out : out std_logic_vector( 72-1 downto 0 );
    ram_1_out : out std_logic_vector( 72-1 downto 0 );
    ram_2_out : out std_logic_vector( 72-1 downto 0 );
    ram_3_out : out std_logic_vector( 72-1 downto 0 );
    ram_4_out : out std_logic_vector( 72-1 downto 0 );
    valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_memory_subsystem;
architecture structural of mh_kernel_memory_subsystem is 
  signal line_out_ram_0_y_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 72-1 downto 0 );
  signal clk_net : std_logic;
  signal line_out_ram_4_y_net : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_2_y_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_3_y_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal remove_offset_mux_read_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 9-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal remove_offset_mux_y_net : std_logic_vector( 9-1 downto 0 );
  signal ce_net : std_logic;
  signal line_out_ram_1_y_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 9-1 downto 0 );
  signal line_out_ram_1_y_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_4_y_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal write_constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal read_constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_doutb_net : std_logic_vector( 72-1 downto 0 );
begin
  ram_0_out <= dual_port_ram_0_douta_net;
  ram_1_out <= dual_port_ram_1_douta_net;
  ram_2_out <= dual_port_ram_2_douta_net;
  ram_3_out <= dual_port_ram_3_douta_net;
  ram_4_out <= dual_port_ram_4_douta_net;
  valid <= convert_to_bool_dout_net;
  remove_offset_mux_y_net <= read_address;
  remove_offset_mux_read_delay_q_net <= read_enable;
  delay_2_q_net <= write_address;
  delay_3_q_net <= write_data_to_ram_sel;
  delay_0_q_net <= data_to_write;
  delay_1_q_net <= write_enable;
  clk_net <= clk_1;
  ce_net <= ce_1;
  ram_selector_0 : entity xil_defaultlib.mh_ram_selector_0 
  port map (
    data_in => delay_2_q_net,
    ram_select => delay_3_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_ram_0 => line_out_ram_0_y_net_x0,
    out_ram_1 => line_out_ram_1_y_net_x0,
    out_ram_2 => line_out_ram_2_y_net_x0,
    out_ram_3 => line_out_ram_3_y_net,
    out_ram_4 => line_out_ram_4_y_net
  );
  ram_selector_1 : entity xil_defaultlib.mh_ram_selector_1 
  port map (
    data_in => delay_0_q_net,
    ram_select => delay_3_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_ram_0 => line_out_ram_0_y_net,
    out_ram_1 => line_out_ram_1_y_net,
    out_ram_2 => line_out_ram_2_y_net,
    out_ram_3 => line_out_ram_3_y_net_x0,
    out_ram_4 => line_out_ram_4_y_net_x0
  );
  ram_selector_2 : entity xil_defaultlib.mh_ram_selector_2_x0 
  port map (
    data_in => delay_1_q_net,
    ram_select => delay_3_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_ram_0 => line_out_ram_0_y_net_x1,
    out_ram_1 => line_out_ram_1_y_net_x1,
    out_ram_2 => line_out_ram_2_y_net_x1,
    out_ram_3 => line_out_ram_3_y_net_x1,
    out_ram_4 => line_out_ram_4_y_net_x1
  );
  convert_to_bool : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => remove_offset_mux_read_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_to_bool_dout_net
  );
  dual_port_ram_0 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 9,
    addr_width_b => 9,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 36000,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_mux_y_net,
    dina => line_out_ram_0_y_net,
    wea => read_constant_op_net,
    addrb => line_out_ram_0_y_net_x0,
    dinb => line_out_ram_0_y_net,
    web => write_constant_op_net,
    ena => remove_offset_mux_read_delay_q_net,
    enb => line_out_ram_0_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 9,
    addr_width_b => 9,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 36000,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_mux_y_net,
    dina => line_out_ram_1_y_net,
    wea => read_constant_op_net,
    addrb => line_out_ram_1_y_net_x0,
    dinb => line_out_ram_1_y_net,
    web => write_constant_op_net,
    ena => remove_offset_mux_read_delay_q_net,
    enb => line_out_ram_1_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  dual_port_ram_2 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 9,
    addr_width_b => 9,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 36000,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_mux_y_net,
    dina => line_out_ram_2_y_net,
    wea => read_constant_op_net,
    addrb => line_out_ram_2_y_net_x0,
    dinb => line_out_ram_2_y_net,
    web => write_constant_op_net,
    ena => remove_offset_mux_read_delay_q_net,
    enb => line_out_ram_2_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_2_douta_net,
    doutb => dual_port_ram_2_doutb_net
  );
  dual_port_ram_3 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 9,
    addr_width_b => 9,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 36000,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_mux_y_net,
    dina => line_out_ram_3_y_net_x0,
    wea => read_constant_op_net,
    addrb => line_out_ram_3_y_net,
    dinb => line_out_ram_3_y_net_x0,
    web => write_constant_op_net,
    ena => remove_offset_mux_read_delay_q_net,
    enb => line_out_ram_3_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_3_douta_net,
    doutb => dual_port_ram_3_doutb_net
  );
  dual_port_ram_4 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 9,
    addr_width_b => 9,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 36000,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_mux_y_net,
    dina => line_out_ram_4_y_net_x0,
    wea => read_constant_op_net,
    addrb => line_out_ram_4_y_net,
    dinb => line_out_ram_4_y_net_x0,
    web => write_constant_op_net,
    ena => remove_offset_mux_read_delay_q_net,
    enb => line_out_ram_4_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_4_douta_net,
    doutb => dual_port_ram_4_doutb_net
  );
  read_constant : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => read_constant_op_net
  );
  write_constant : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => write_constant_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Memory Sync
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_memory_sync is
  port (
    frame_memory_full : in std_logic_vector( 1-1 downto 0 );
    kernel_memory_full : in std_logic_vector( 1-1 downto 0 );
    new_frame : in std_logic_vector( 1-1 downto 0 );
    reset : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    frame_memory_address : out std_logic_vector( 17-1 downto 0 );
    frame_read_enable : out std_logic_vector( 1-1 downto 0 );
    kernel_memory_address : out std_logic_vector( 9-1 downto 0 );
    kernel_read_enable : out std_logic_vector( 1-1 downto 0 )
  );
end mh_memory_sync;
architecture structural of mh_memory_sync is 
  signal hold_up_read_out_frame_op_net : std_logic_vector( 1-1 downto 0 );
  signal remove_offset_frame_memory_address_delay_q_net : std_logic_vector( 17-1 downto 0 );
  signal remove_offset_frame_read_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal subtrack_frame_memory_address_delay_q_net : std_logic_vector( 17-1 downto 0 );
  signal subtrack_frame_read_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal subtrack_kernel_read_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal remove_offset_original_delay_and_cast_dout_net : std_logic_vector( 9-1 downto 0 );
  signal remove_offset_subtracked_delay_and_cast_dout_net : std_logic_vector( 9-1 downto 0 );
  signal subtrack_offset_s_net : std_logic_vector( 11-1 downto 0 );
  signal remove_offset_kernel_read_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal remove_offset_frame_memory_address_delay1_q_net : std_logic_vector( 17-1 downto 0 );
  signal remove_offset_mux_y_net : std_logic_vector( 9-1 downto 0 );
  signal memory_full_delay_2_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal memory_full_delay_1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal add_frame_memory_address_delay_q_net : std_logic_vector( 17-1 downto 0 );
  signal count_to_max_frame_memory_op_net : std_logic_vector( 17-1 downto 0 );
  signal memory_full_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal remove_offset_frame_read_enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_frame_read_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal frame_counter_all_on_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal remove_offset_mux_read_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant1_op_net_x0 : std_logic_vector( 2-1 downto 0 );
  signal check_once1_y_net : std_logic_vector( 1-1 downto 0 );
  signal kernel_offset_op_net : std_logic_vector( 9-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 8-1 downto 0 );
  signal kernel_count_full_op_net : std_logic_vector( 9-1 downto 0 );
  signal check_to_remove_offset_op_net : std_logic_vector( 1-1 downto 0 );
  signal subtrack_delay_q_net : std_logic_vector( 10-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 9-1 downto 0 );
  signal add_offset_s_net : std_logic_vector( 10-1 downto 0 );
  signal check_if_2_frame_sync_op_net : std_logic_vector( 1-1 downto 0 );
  signal check_if_at_reset_point_op_net : std_logic_vector( 1-1 downto 0 );
  signal count_to_3_op_net : std_logic_vector( 2-1 downto 0 );
  signal add_kernel_read_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal turn_on_generator_dout_net : std_logic_vector( 1-1 downto 0 );
  signal check_last_address1_op_net : std_logic_vector( 1-1 downto 0 );
  signal kernel_count_op_net : std_logic_vector( 7-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 9-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_circular_buffer_state_update_q_net : std_logic_vector( 1-1 downto 0 );
  signal count_positive_y_net : std_logic_vector( 1-1 downto 0 );
  signal enable_frame_counter_y_net : std_logic_vector( 1-1 downto 0 );
begin
  frame_memory_address <= remove_offset_frame_memory_address_delay1_q_net;
  frame_read_enable <= remove_offset_frame_read_enable_delay1_q_net;
  kernel_memory_address <= remove_offset_mux_y_net;
  kernel_read_enable <= remove_offset_mux_read_delay_q_net;
  memory_full_delay_1_q_net_x0 <= frame_memory_full;
  memory_full_delay_1_q_net <= kernel_memory_full;
  memory_full_delay_2_q_net <= new_frame;
  constant1_op_net <= reset;
  clk_net <= clk_1;
  ce_net <= ce_1;
  add_frame_memory_address_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 17
  )
  port map (
    en => '1',
    rst => '0',
    d => count_to_max_frame_memory_op_net,
    clk => clk_net,
    ce => ce_net,
    q => add_frame_memory_address_delay_q_net
  );
  add_frame_read_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => frame_counter_all_on_y_net,
    clk => clk_net,
    ce => ce_net,
    q => add_frame_read_enable_delay_q_net
  );
  add_kernel_read_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => turn_on_generator_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => add_kernel_read_enable_delay_q_net
  );
  add_offset : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 9,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 9,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 10,
    core_name0 => "mh_c_addsub_v12_0_i9",
    extra_registers => 0,
    full_s_arith => 1,
    full_s_width => 10,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 10
  )
  port map (
    clr => '0',
    en => "1",
    a => kernel_count_full_op_net,
    b => kernel_offset_op_net,
    clk => clk_net,
    ce => ce_net,
    s => add_offset_s_net
  );
  check_if_at_reset_point : entity xil_defaultlib.sysgen_relational_2751815a1d 
  port map (
    clr => '0',
    a => constant5_op_net,
    b => kernel_count_op_net,
    clk => clk_net,
    ce => ce_net,
    op => check_if_at_reset_point_op_net
  );
  check_last_address1 : entity xil_defaultlib.sysgen_relational_7e7f05af27 
  port map (
    clr => '0',
    a => count_to_max_frame_memory_op_net,
    b => constant2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => check_last_address1_op_net
  );
  check_once1 : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => delay1_q_net,
    d1 => check_last_address1_op_net,
    clk => clk_net,
    ce => ce_net,
    y => check_once1_y_net
  );
  check_if_2_frame_sync : entity xil_defaultlib.sysgen_relational_7e2637e235 
  port map (
    clr => '0',
    a => constant1_op_net_x0,
    b => count_to_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => check_if_2_frame_sync_op_net
  );
  check_to_remove_offset : entity xil_defaultlib.sysgen_relational_affb8e2e51 
  port map (
    clr => '0',
    a => subtrack_delay_q_net,
    b => constant3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => check_to_remove_offset_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_9d2d62a34e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net_x0
  );
  constant2 : entity xil_defaultlib.sysgen_constant_abbf85fae7 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_d8cf2ae02b 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_4a0587bd7f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_44931d96aa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  count_positive : entity xil_defaultlib.sysgen_logical_5b21a0b250 
  port map (
    clr => '0',
    d0 => logical_y_net,
    d1 => constant1_op_net,
    clk => clk_net,
    ce => ce_net,
    y => count_positive_y_net
  );
  count_to_3 : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 2,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i1",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => check_if_at_reset_point_op_net,
    en => turn_on_generator_dout_net,
    clk => clk_net,
    ce => ce_net,
    op => count_to_3_op_net
  );
  count_to_max_frame_memory : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 8163,
    cnt_31_16 => 1,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i18",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 17
  )
  port map (
    rst => "0",
    clr => '0',
    en => frame_counter_all_on_y_net,
    clk => clk_net,
    ce => ce_net,
    op => count_to_max_frame_memory_op_net
  );
  delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => frame_counter_all_on_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  enable_circular_buffer_state_update : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => check_once1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => enable_circular_buffer_state_update_q_net
  );
  enable_frame_counter : entity xil_defaultlib.sysgen_logical_b4b46f5c45 
  port map (
    clr => '0',
    d0 => logical_y_net,
    d1 => constant1_op_net,
    d2 => check_once1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => enable_frame_counter_y_net
  );
  frame_counter_all_on : entity xil_defaultlib.sysgen_logical_f780ce33fa 
  port map (
    clr => '0',
    d0 => check_if_2_frame_sync_op_net,
    d1 => turn_on_generator_dout_net,
    clk => clk_net,
    ce => ce_net,
    y => frame_counter_all_on_y_net
  );
  hold_up_read_out_frame : entity xil_defaultlib.sysgen_counter_1070c7a3c7 
  port map (
    clr => '0',
    up => count_positive_y_net,
    en => enable_frame_counter_y_net,
    clk => clk_net,
    ce => ce_net,
    op => hold_up_read_out_frame_op_net
  );
  kernel_count : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 99,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i0",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    rst => "0",
    clr => '0',
    en => turn_on_generator_dout_net,
    clk => clk_net,
    ce => ce_net,
    op => kernel_count_op_net
  );
  kernel_count_full : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 499,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i10",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => turn_on_generator_dout_net,
    clk => clk_net,
    ce => ce_net,
    op => kernel_count_full_op_net
  );
  kernel_offset : entity xil_defaultlib.mh_xlcounter_limit 
  generic map (
    cnt_15_0 => 100,
    cnt_31_16 => 0,
    cnt_47_32 => 0,
    cnt_63_48 => 0,
    core_name0 => "mh_c_counter_binary_v12_0_i19",
    count_limited => 1,
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    rst => "0",
    clr => '0',
    en => enable_circular_buffer_state_update_q_net,
    clk => clk_net,
    ce => ce_net,
    op => kernel_offset_op_net
  );
  logical : entity xil_defaultlib.sysgen_logical_8d46e13166 
  port map (
    clr => '0',
    d0 => memory_full_delay_1_q_net_x0,
    d1 => memory_full_delay_1_q_net,
    d2 => memory_full_delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  remove_offset_frame_memory_address_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 17
  )
  port map (
    en => '1',
    rst => '0',
    d => subtrack_frame_memory_address_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => remove_offset_frame_memory_address_delay_q_net
  );
  remove_offset_frame_memory_address_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 17
  )
  port map (
    en => '1',
    rst => '0',
    d => remove_offset_frame_memory_address_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => remove_offset_frame_memory_address_delay1_q_net
  );
  remove_offset_frame_read_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => subtrack_frame_read_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => remove_offset_frame_read_enable_delay_q_net
  );
  remove_offset_frame_read_enable_delay1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => remove_offset_frame_read_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => remove_offset_frame_read_enable_delay1_q_net
  );
  remove_offset_kernel_read_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => subtrack_kernel_read_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => remove_offset_kernel_read_delay_q_net
  );
  remove_offset_mux : entity xil_defaultlib.sysgen_mux_044d346e3b 
  port map (
    clr => '0',
    sel => check_to_remove_offset_op_net,
    d0 => remove_offset_subtracked_delay_and_cast_dout_net,
    d1 => remove_offset_original_delay_and_cast_dout_net,
    clk => clk_net,
    ce => ce_net,
    y => remove_offset_mux_y_net
  );
  remove_offset_mux_read_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => remove_offset_kernel_read_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => remove_offset_mux_read_delay_q_net
  );
  remove_offset_original_delay_and_cast : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 0,
    din_width => 11,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 9,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => subtrack_offset_s_net,
    clk => clk_net,
    ce => ce_net,
    dout => remove_offset_original_delay_and_cast_dout_net
  );
  remove_offset_subtracked_delay_and_cast : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 10,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 9,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => subtrack_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    dout => remove_offset_subtracked_delay_and_cast_dout_net
  );
  subtrack_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 10
  )
  port map (
    en => '1',
    rst => '0',
    d => add_offset_s_net,
    clk => clk_net,
    ce => ce_net,
    q => subtrack_delay_q_net
  );
  subtrack_frame_memory_address_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 17
  )
  port map (
    en => '1',
    rst => '0',
    d => add_frame_memory_address_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => subtrack_frame_memory_address_delay_q_net
  );
  subtrack_frame_read_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => add_frame_read_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => subtrack_frame_read_enable_delay_q_net
  );
  subtrack_kernel_read_enable_delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => add_kernel_read_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => subtrack_kernel_read_enable_delay_q_net
  );
  subtrack_offset : entity xil_defaultlib.mh_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 10,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 9,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 11,
    core_name0 => "mh_c_addsub_v12_0_i10",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 11,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 0,
    s_width => 11
  )
  port map (
    clr => '0',
    en => "1",
    a => add_offset_s_net,
    b => constant4_op_net,
    clk => clk_net,
    ce => ce_net,
    s => subtrack_offset_s_net
  );
  turn_on_generator : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => hold_up_read_out_frame_op_net,
    clk => clk_net,
    ce => ce_net,
    dout => turn_on_generator_dout_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Memory Sync Delay Frame Write
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_memory_sync_delay_frame_write is
  port (
    data_out_72_bits : in std_logic_vector( 72-1 downto 0 );
    data_out_ready : in std_logic_vector( 1-1 downto 0 );
    data_address_out : in std_logic_vector( 17-1 downto 0 );
    ram_bloack_sel_out : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_to_write : out std_logic_vector( 72-1 downto 0 );
    write_enable : out std_logic_vector( 1-1 downto 0 );
    write_address : out std_logic_vector( 17-1 downto 0 );
    write_data_to_ram_sel : out std_logic_vector( 3-1 downto 0 )
  );
end mh_memory_sync_delay_frame_write;
architecture structural of mh_memory_sync_delay_frame_write is 
  signal final_add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal add_ram_sel_delay_1_q_net : std_logic_vector( 3-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal final_add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_offset_with_line_count_s_net : std_logic_vector( 17-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 17-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
begin
  data_to_write <= delay_0_q_net;
  write_enable <= delay_1_q_net;
  write_address <= delay_2_q_net;
  write_data_to_ram_sel <= delay_3_q_net;
  final_add_data_out_delay_q_net <= data_out_72_bits;
  final_add_enable_delay_q_net <= data_out_ready;
  add_offset_with_line_count_s_net <= data_address_out;
  add_ram_sel_delay_1_q_net <= ram_bloack_sel_out;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 600,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => final_add_data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_0_q_net
  );
  delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 600,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => final_add_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_1_q_net
  );
  delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 600,
    reg_retiming => 0,
    reset => 0,
    width => 17
  )
  port map (
    en => '1',
    rst => '0',
    d => add_offset_with_line_count_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_2_q_net
  );
  delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 600,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => add_ram_sel_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_3_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Memory Sync Delay Frame Write1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_memory_sync_delay_frame_write1 is
  port (
    data_out_72_bits : in std_logic_vector( 72-1 downto 0 );
    data_out_ready : in std_logic_vector( 1-1 downto 0 );
    data_address_out : in std_logic_vector( 9-1 downto 0 );
    ram_bloack_sel_out : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_to_write : out std_logic_vector( 72-1 downto 0 );
    write_enable : out std_logic_vector( 1-1 downto 0 );
    write_address : out std_logic_vector( 9-1 downto 0 );
    write_data_to_ram_sel : out std_logic_vector( 3-1 downto 0 )
  );
end mh_memory_sync_delay_frame_write1;
architecture structural of mh_memory_sync_delay_frame_write1 is 
  signal final_add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal final_add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal ce_net : std_logic;
  signal data_out_delay_q_net : std_logic_vector( 9-1 downto 0 );
  signal add_ram_sel_delay_1_q_net : std_logic_vector( 3-1 downto 0 );
  signal clk_net : std_logic;
begin
  data_to_write <= delay_0_q_net;
  write_enable <= delay_1_q_net;
  write_address <= delay_2_q_net;
  write_data_to_ram_sel <= delay_3_q_net;
  final_add_data_out_delay_q_net <= data_out_72_bits;
  final_add_enable_delay_q_net <= data_out_ready;
  data_out_delay_q_net <= data_address_out;
  add_ram_sel_delay_1_q_net <= ram_bloack_sel_out;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay_0 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 400,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => final_add_data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_0_q_net
  );
  delay_1 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 400,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => final_add_enable_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_1_q_net
  );
  delay_2 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 400,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => data_out_delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_2_q_net
  );
  delay_3 : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 400,
    reg_retiming => 0,
    reset => 0,
    width => 3
  )
  port map (
    en => '1',
    rst => '0',
    d => add_ram_sel_delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_3_q_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Scanline Memory Subsystem/RAM Selector 0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_ram_selector_0_x0 is
  port (
    data_in : in std_logic_vector( 17-1 downto 0 );
    ram_select : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_ram_0 : out std_logic_vector( 17-1 downto 0 );
    out_ram_1 : out std_logic_vector( 17-1 downto 0 );
    out_ram_2 : out std_logic_vector( 17-1 downto 0 );
    out_ram_3 : out std_logic_vector( 17-1 downto 0 );
    out_ram_4 : out std_logic_vector( 17-1 downto 0 )
  );
end mh_ram_selector_0_x0;
architecture structural of mh_ram_selector_0_x0 is 
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 17-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 17-1 downto 0 );
  signal line_out_ram_4_y_net : std_logic_vector( 17-1 downto 0 );
  signal ce_net : std_logic;
  signal line_out_ram_1_y_net : std_logic_vector( 17-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 17-1 downto 0 );
  signal sel_value_ram_1_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_2_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_0_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_4_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_3_op_net : std_logic_vector( 3-1 downto 0 );
begin
  out_ram_0 <= line_out_ram_0_y_net;
  out_ram_1 <= line_out_ram_1_y_net;
  out_ram_2 <= line_out_ram_2_y_net;
  out_ram_3 <= line_out_ram_3_y_net;
  out_ram_4 <= line_out_ram_4_y_net;
  delay_2_q_net <= data_in;
  delay_3_q_net <= ram_select;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 17
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  line_out_ram_0 : entity xil_defaultlib.sysgen_mux_f38fc9b1d2 
  port map (
    clr => '0',
    sel => sel_ram_0_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_0_y_net
  );
  line_out_ram_1 : entity xil_defaultlib.sysgen_mux_f38fc9b1d2 
  port map (
    clr => '0',
    sel => sel_ram_1_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_1_y_net
  );
  line_out_ram_2 : entity xil_defaultlib.sysgen_mux_f38fc9b1d2 
  port map (
    clr => '0',
    sel => sel_ram_2_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_2_y_net
  );
  line_out_ram_3 : entity xil_defaultlib.sysgen_mux_f38fc9b1d2 
  port map (
    clr => '0',
    sel => sel_ram_3_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_3_y_net
  );
  line_out_ram_4 : entity xil_defaultlib.sysgen_mux_f38fc9b1d2 
  port map (
    clr => '0',
    sel => sel_ram_4_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_4_y_net
  );
  sel_ram_0 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_0_op_net
  );
  sel_ram_1 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_1_op_net
  );
  sel_ram_2 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_2_op_net
  );
  sel_ram_3 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_3_op_net
  );
  sel_ram_4 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_4_op_net
  );
  sel_value_ram_0 : entity xil_defaultlib.sysgen_constant_28e1aa0294 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_0_op_net
  );
  sel_value_ram_1 : entity xil_defaultlib.sysgen_constant_031f960172 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_1_op_net
  );
  sel_value_ram_2 : entity xil_defaultlib.sysgen_constant_15681d4665 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_2_op_net
  );
  sel_value_ram_3 : entity xil_defaultlib.sysgen_constant_c571582d8a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_3_op_net
  );
  sel_value_ram_4 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_4_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Scanline Memory Subsystem/RAM Selector 1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_ram_selector_1_x0 is
  port (
    data_in : in std_logic_vector( 72-1 downto 0 );
    ram_select : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_ram_0 : out std_logic_vector( 72-1 downto 0 );
    out_ram_1 : out std_logic_vector( 72-1 downto 0 );
    out_ram_2 : out std_logic_vector( 72-1 downto 0 );
    out_ram_3 : out std_logic_vector( 72-1 downto 0 );
    out_ram_4 : out std_logic_vector( 72-1 downto 0 )
  );
end mh_ram_selector_1_x0;
architecture structural of mh_ram_selector_1_x0 is 
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_4_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_1_y_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 72-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal sel_ram_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_0_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_1_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_2_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_3_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_4_op_net : std_logic_vector( 3-1 downto 0 );
begin
  out_ram_0 <= line_out_ram_0_y_net;
  out_ram_1 <= line_out_ram_1_y_net;
  out_ram_2 <= line_out_ram_2_y_net;
  out_ram_3 <= line_out_ram_3_y_net;
  out_ram_4 <= line_out_ram_4_y_net;
  delay_0_q_net <= data_in;
  delay_3_q_net <= ram_select;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 72
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  line_out_ram_0 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_0_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_0_y_net
  );
  line_out_ram_1 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_1_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_1_y_net
  );
  line_out_ram_2 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_2_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_2_y_net
  );
  line_out_ram_3 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_3_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_3_y_net
  );
  line_out_ram_4 : entity xil_defaultlib.sysgen_mux_decbbe2618 
  port map (
    clr => '0',
    sel => sel_ram_4_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_4_y_net
  );
  sel_ram_0 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_0_op_net
  );
  sel_ram_1 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_1_op_net
  );
  sel_ram_2 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_2_op_net
  );
  sel_ram_3 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_3_op_net
  );
  sel_ram_4 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_4_op_net
  );
  sel_value_ram_0 : entity xil_defaultlib.sysgen_constant_28e1aa0294 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_0_op_net
  );
  sel_value_ram_1 : entity xil_defaultlib.sysgen_constant_031f960172 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_1_op_net
  );
  sel_value_ram_2 : entity xil_defaultlib.sysgen_constant_15681d4665 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_2_op_net
  );
  sel_value_ram_3 : entity xil_defaultlib.sysgen_constant_c571582d8a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_3_op_net
  );
  sel_value_ram_4 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_4_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Scanline Memory Subsystem/RAM Selector 2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_ram_selector_2 is
  port (
    data_in : in std_logic_vector( 1-1 downto 0 );
    ram_select : in std_logic_vector( 3-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_ram_0 : out std_logic_vector( 1-1 downto 0 );
    out_ram_1 : out std_logic_vector( 1-1 downto 0 );
    out_ram_2 : out std_logic_vector( 1-1 downto 0 );
    out_ram_3 : out std_logic_vector( 1-1 downto 0 );
    out_ram_4 : out std_logic_vector( 1-1 downto 0 )
  );
end mh_ram_selector_2;
architecture structural of mh_ram_selector_2 is 
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal line_out_ram_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_1_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_4_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_2_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_3_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_1_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_3_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_ram_0_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_ram_2_op_net : std_logic_vector( 1-1 downto 0 );
  signal sel_value_ram_0_op_net : std_logic_vector( 3-1 downto 0 );
  signal sel_value_ram_4_op_net : std_logic_vector( 3-1 downto 0 );
begin
  out_ram_0 <= line_out_ram_0_y_net;
  out_ram_1 <= line_out_ram_1_y_net;
  out_ram_2 <= line_out_ram_2_y_net;
  out_ram_3 <= line_out_ram_3_y_net;
  out_ram_4 <= line_out_ram_4_y_net;
  delay_1_q_net <= data_in;
  delay_3_q_net <= ram_select;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.mh_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay_1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  line_out_ram_0 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_0_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_0_y_net
  );
  line_out_ram_1 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_1_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_1_y_net
  );
  line_out_ram_2 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_2_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_2_y_net
  );
  line_out_ram_3 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_3_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_3_y_net
  );
  line_out_ram_4 : entity xil_defaultlib.sysgen_mux_41e92c8c2c 
  port map (
    clr => '0',
    sel => sel_ram_4_op_net,
    d0 => constant1_op_net,
    d1 => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    y => line_out_ram_4_y_net
  );
  sel_ram_0 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_0_op_net
  );
  sel_ram_1 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_1_op_net
  );
  sel_ram_2 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_2_op_net
  );
  sel_ram_3 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_3_op_net
  );
  sel_ram_4 : entity xil_defaultlib.sysgen_relational_4ad15b3c66 
  port map (
    clr => '0',
    a => delay_3_q_net,
    b => sel_value_ram_4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => sel_ram_4_op_net
  );
  sel_value_ram_0 : entity xil_defaultlib.sysgen_constant_28e1aa0294 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_0_op_net
  );
  sel_value_ram_1 : entity xil_defaultlib.sysgen_constant_031f960172 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_1_op_net
  );
  sel_value_ram_2 : entity xil_defaultlib.sysgen_constant_15681d4665 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_2_op_net
  );
  sel_value_ram_3 : entity xil_defaultlib.sysgen_constant_c571582d8a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_3_op_net
  );
  sel_value_ram_4 : entity xil_defaultlib.sysgen_constant_348be6236f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => sel_value_ram_4_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Scanline Memory Subsystem
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_scanline_memory_subsystem is
  port (
    read_address : in std_logic_vector( 17-1 downto 0 );
    read_enable : in std_logic_vector( 1-1 downto 0 );
    write_address : in std_logic_vector( 17-1 downto 0 );
    write_data_to_ram_sel : in std_logic_vector( 3-1 downto 0 );
    data_to_write : in std_logic_vector( 72-1 downto 0 );
    write_enable : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ram_0_out : out std_logic_vector( 72-1 downto 0 );
    ram_1_out : out std_logic_vector( 72-1 downto 0 );
    ram_2_out : out std_logic_vector( 72-1 downto 0 );
    ram_3_out : out std_logic_vector( 72-1 downto 0 );
    ram_4_out : out std_logic_vector( 72-1 downto 0 );
    valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_scanline_memory_subsystem;
architecture structural of mh_scanline_memory_subsystem is 
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal line_out_ram_1_y_net : std_logic_vector( 17-1 downto 0 );
  signal line_out_ram_2_y_net : std_logic_vector( 17-1 downto 0 );
  signal line_out_ram_3_y_net_x0 : std_logic_vector( 17-1 downto 0 );
  signal line_out_ram_0_y_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal remove_offset_frame_memory_address_delay1_q_net : std_logic_vector( 17-1 downto 0 );
  signal ce_net : std_logic;
  signal line_out_ram_0_y_net : std_logic_vector( 17-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_4_y_net_x0 : std_logic_vector( 17-1 downto 0 );
  signal line_out_ram_1_y_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_2_y_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_3_y_net_x1 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal remove_offset_frame_read_enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 17-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal read_constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal line_out_ram_4_y_net_x1 : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal write_constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal line_out_ram_0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_3_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_doutb_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_doutb_net : std_logic_vector( 72-1 downto 0 );
begin
  ram_0_out <= dual_port_ram_0_douta_net;
  ram_1_out <= dual_port_ram_1_douta_net;
  ram_2_out <= dual_port_ram_2_douta_net;
  ram_3_out <= dual_port_ram_3_douta_net;
  ram_4_out <= dual_port_ram_4_douta_net;
  valid <= convert_to_bool_dout_net;
  remove_offset_frame_memory_address_delay1_q_net <= read_address;
  remove_offset_frame_read_enable_delay1_q_net <= read_enable;
  delay_2_q_net <= write_address;
  delay_3_q_net <= write_data_to_ram_sel;
  delay_0_q_net <= data_to_write;
  delay_1_q_net <= write_enable;
  clk_net <= clk_1;
  ce_net <= ce_1;
  ram_selector_0 : entity xil_defaultlib.mh_ram_selector_0_x0 
  port map (
    data_in => delay_2_q_net,
    ram_select => delay_3_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_ram_0 => line_out_ram_0_y_net,
    out_ram_1 => line_out_ram_1_y_net,
    out_ram_2 => line_out_ram_2_y_net,
    out_ram_3 => line_out_ram_3_y_net_x0,
    out_ram_4 => line_out_ram_4_y_net_x0
  );
  ram_selector_1 : entity xil_defaultlib.mh_ram_selector_1_x0 
  port map (
    data_in => delay_0_q_net,
    ram_select => delay_3_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_ram_0 => line_out_ram_0_y_net_x0,
    out_ram_1 => line_out_ram_1_y_net_x0,
    out_ram_2 => line_out_ram_2_y_net_x0,
    out_ram_3 => line_out_ram_3_y_net_x1,
    out_ram_4 => line_out_ram_4_y_net_x1
  );
  ram_selector_2 : entity xil_defaultlib.mh_ram_selector_2 
  port map (
    data_in => delay_1_q_net,
    ram_select => delay_3_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_ram_0 => line_out_ram_0_y_net_x1,
    out_ram_1 => line_out_ram_1_y_net_x1,
    out_ram_2 => line_out_ram_2_y_net_x1,
    out_ram_3 => line_out_ram_3_y_net,
    out_ram_4 => line_out_ram_4_y_net
  );
  convert_to_bool : entity xil_defaultlib.mh_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => remove_offset_frame_read_enable_delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_to_bool_dout_net
  );
  dual_port_ram_0 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 17,
    addr_width_b => 17,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 5306400,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_frame_memory_address_delay1_q_net,
    dina => line_out_ram_0_y_net_x0,
    wea => read_constant_op_net,
    addrb => line_out_ram_0_y_net,
    dinb => line_out_ram_0_y_net_x0,
    web => write_constant_op_net,
    ena => remove_offset_frame_read_enable_delay1_q_net,
    enb => line_out_ram_0_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 17,
    addr_width_b => 17,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 5306400,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_frame_memory_address_delay1_q_net,
    dina => line_out_ram_1_y_net_x0,
    wea => read_constant_op_net,
    addrb => line_out_ram_1_y_net,
    dinb => line_out_ram_1_y_net_x0,
    web => write_constant_op_net,
    ena => remove_offset_frame_read_enable_delay1_q_net,
    enb => line_out_ram_1_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  dual_port_ram_2 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 17,
    addr_width_b => 17,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 5306400,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_frame_memory_address_delay1_q_net,
    dina => line_out_ram_2_y_net_x0,
    wea => read_constant_op_net,
    addrb => line_out_ram_2_y_net,
    dinb => line_out_ram_2_y_net_x0,
    web => write_constant_op_net,
    ena => remove_offset_frame_read_enable_delay1_q_net,
    enb => line_out_ram_2_y_net_x1,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_2_douta_net,
    doutb => dual_port_ram_2_doutb_net
  );
  dual_port_ram_3 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 17,
    addr_width_b => 17,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 5306400,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_frame_memory_address_delay1_q_net,
    dina => line_out_ram_3_y_net_x1,
    wea => read_constant_op_net,
    addrb => line_out_ram_3_y_net_x0,
    dinb => line_out_ram_3_y_net_x1,
    web => write_constant_op_net,
    ena => remove_offset_frame_read_enable_delay1_q_net,
    enb => line_out_ram_3_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_3_douta_net,
    doutb => dual_port_ram_3_doutb_net
  );
  dual_port_ram_4 : entity xil_defaultlib.mh_xltdpram 
  generic map (
    addr_width_a => 17,
    addr_width_b => 17,
    data_width_a => 72,
    data_width_b => 72,
    latency => 1,
    mem_size => 5306400,
    mem_type => "ultra",
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    rsta => "0",
    rstb => "0",
    addra => remove_offset_frame_memory_address_delay1_q_net,
    dina => line_out_ram_4_y_net_x1,
    wea => read_constant_op_net,
    addrb => line_out_ram_4_y_net_x0,
    dinb => line_out_ram_4_y_net_x1,
    web => write_constant_op_net,
    ena => remove_offset_frame_read_enable_delay1_q_net,
    enb => line_out_ram_4_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_4_douta_net,
    doutb => dual_port_ram_4_doutb_net
  );
  read_constant : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => read_constant_op_net
  );
  write_constant : entity xil_defaultlib.sysgen_constant_3dd30f50e6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => write_constant_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_memory_manager is
  port (
    x12_bit_spectrual_bin_in : in std_logic_vector( 12-1 downto 0 );
    enable_in_spectrual : in std_logic_vector( 1-1 downto 0 );
    x18_bit_kernel_data_in : in std_logic_vector( 18-1 downto 0 );
    enable_in_kernel : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    spectrual_ram_0_out : out std_logic_vector( 72-1 downto 0 );
    spectrual_ram_1_out : out std_logic_vector( 72-1 downto 0 );
    spectrual_ram_2_out : out std_logic_vector( 72-1 downto 0 );
    spectrual_ram_3_out : out std_logic_vector( 72-1 downto 0 );
    spectrual_ram_4_out : out std_logic_vector( 72-1 downto 0 );
    spectrual_valid : out std_logic_vector( 1-1 downto 0 );
    kernel_ram_0_out1 : out std_logic_vector( 72-1 downto 0 );
    kernel_ram_1_out1 : out std_logic_vector( 72-1 downto 0 );
    kernel_ram_2_out1 : out std_logic_vector( 72-1 downto 0 );
    kernel_ram_3_out1 : out std_logic_vector( 72-1 downto 0 );
    kernel_ram_4_out1 : out std_logic_vector( 72-1 downto 0 );
    kernel_valid : out std_logic_vector( 1-1 downto 0 )
  );
end mh_memory_manager;
architecture structural of mh_memory_manager is 
  signal dual_port_ram_0_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_1_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal remove_offset_frame_memory_address_delay1_q_net : std_logic_vector( 17-1 downto 0 );
  signal add_offset_with_line_count_s_net : std_logic_vector( 17-1 downto 0 );
  signal delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal memory_full_delay_2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal final_add_data_out_delay_q_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal remove_offset_frame_read_enable_delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_18_bit_net : std_logic_vector( 18-1 downto 0 );
  signal final_add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_ram_sel_delay_1_q_net : std_logic_vector( 3-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal write_enable_12_bit_net : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net_x0 : std_logic_vector( 17-1 downto 0 );
  signal delay_3_q_net : std_logic_vector( 3-1 downto 0 );
  signal convert_to_bool_dout_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal memory_full_delay_1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_2_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay_0_q_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal ce_net : std_logic;
  signal data_out_delay_q_net : std_logic_vector( 9-1 downto 0 );
  signal final_add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal memory_full_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal remove_offset_mux_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay_0_q_net : std_logic_vector( 72-1 downto 0 );
  signal delay_1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay_3_q_net_x0 : std_logic_vector( 3-1 downto 0 );
  signal remove_offset_mux_read_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_enable_18_bit_net : std_logic_vector( 1-1 downto 0 );
  signal add_ram_sel_delay_1_q_net_x0 : std_logic_vector( 3-1 downto 0 );
  signal final_add_enable_delay_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal data_input_12_bit_net : std_logic_vector( 12-1 downto 0 );
begin
  spectrual_ram_0_out <= dual_port_ram_0_douta_net_x0;
  spectrual_ram_1_out <= dual_port_ram_1_douta_net_x0;
  spectrual_ram_2_out <= dual_port_ram_2_douta_net_x0;
  spectrual_ram_3_out <= dual_port_ram_3_douta_net_x0;
  spectrual_ram_4_out <= dual_port_ram_4_douta_net_x0;
  spectrual_valid <= convert_to_bool_dout_net;
  kernel_ram_0_out1 <= dual_port_ram_0_douta_net;
  kernel_ram_1_out1 <= dual_port_ram_1_douta_net;
  kernel_ram_2_out1 <= dual_port_ram_2_douta_net;
  kernel_ram_3_out1 <= dual_port_ram_3_douta_net;
  kernel_ram_4_out1 <= dual_port_ram_4_douta_net;
  kernel_valid <= convert_to_bool_dout_net_x0;
  data_input_12_bit_net <= x12_bit_spectrual_bin_in;
  write_enable_12_bit_net <= enable_in_spectrual;
  data_in_18_bit_net <= x18_bit_kernel_data_in;
  data_enable_18_bit_net <= enable_in_kernel;
  clk_net <= clk_1;
  ce_net <= ce_1;
  frame_memory_controller : entity xil_defaultlib.mh_frame_memory_controller 
  port map (
    x12_bit_data_in => data_input_12_bit_net,
    enable_in => write_enable_12_bit_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    data_out_72_bits => final_add_data_out_delay_q_net_x0,
    data_out_ready => final_add_enable_delay_q_net_x0,
    data_address_out => add_offset_with_line_count_s_net,
    ram_bloack_sel_out => add_ram_sel_delay_1_q_net_x0,
    memory_is_full => memory_full_delay_1_q_net_x0,
    new_frame_finished => memory_full_delay_2_q_net_x0
  );
  kernel_memory_controller : entity xil_defaultlib.mh_kernel_memory_controller 
  port map (
    x18_bit_data_in => data_in_18_bit_net,
    enable_in => data_enable_18_bit_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    data_out_72_bits => final_add_data_out_delay_q_net,
    data_out_ready => final_add_enable_delay_q_net,
    data_address_out => data_out_delay_q_net,
    ram_block_sel_out => add_ram_sel_delay_1_q_net,
    memory_is_full => memory_full_delay_1_q_net
  );
  kernel_memory_subsystem : entity xil_defaultlib.mh_kernel_memory_subsystem 
  port map (
    read_address => remove_offset_mux_y_net,
    read_enable => remove_offset_mux_read_delay_q_net,
    write_address => delay_2_q_net,
    write_data_to_ram_sel => delay_3_q_net,
    data_to_write => delay_0_q_net,
    write_enable => delay_1_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ram_0_out => dual_port_ram_0_douta_net,
    ram_1_out => dual_port_ram_1_douta_net,
    ram_2_out => dual_port_ram_2_douta_net,
    ram_3_out => dual_port_ram_3_douta_net,
    ram_4_out => dual_port_ram_4_douta_net,
    valid => convert_to_bool_dout_net_x0
  );
  memory_sync : entity xil_defaultlib.mh_memory_sync 
  port map (
    frame_memory_full => memory_full_delay_1_q_net_x0,
    kernel_memory_full => memory_full_delay_1_q_net,
    new_frame => memory_full_delay_2_q_net_x0,
    reset => constant1_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    frame_memory_address => remove_offset_frame_memory_address_delay1_q_net,
    frame_read_enable => remove_offset_frame_read_enable_delay1_q_net,
    kernel_memory_address => remove_offset_mux_y_net,
    kernel_read_enable => remove_offset_mux_read_delay_q_net
  );
  memory_sync_delay_frame_write : entity xil_defaultlib.mh_memory_sync_delay_frame_write 
  port map (
    data_out_72_bits => final_add_data_out_delay_q_net_x0,
    data_out_ready => final_add_enable_delay_q_net_x0,
    data_address_out => add_offset_with_line_count_s_net,
    ram_bloack_sel_out => add_ram_sel_delay_1_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    data_to_write => delay_0_q_net_x0,
    write_enable => delay_1_q_net_x0,
    write_address => delay_2_q_net_x0,
    write_data_to_ram_sel => delay_3_q_net_x0
  );
  memory_sync_delay_frame_write1 : entity xil_defaultlib.mh_memory_sync_delay_frame_write1 
  port map (
    data_out_72_bits => final_add_data_out_delay_q_net,
    data_out_ready => final_add_enable_delay_q_net,
    data_address_out => data_out_delay_q_net,
    ram_bloack_sel_out => add_ram_sel_delay_1_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    data_to_write => delay_0_q_net,
    write_enable => delay_1_q_net,
    write_address => delay_2_q_net,
    write_data_to_ram_sel => delay_3_q_net
  );
  scanline_memory_subsystem : entity xil_defaultlib.mh_scanline_memory_subsystem 
  port map (
    read_address => remove_offset_frame_memory_address_delay1_q_net,
    read_enable => remove_offset_frame_read_enable_delay1_q_net,
    write_address => delay_2_q_net_x0,
    write_data_to_ram_sel => delay_3_q_net_x0,
    data_to_write => delay_0_q_net_x0,
    write_enable => delay_1_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ram_0_out => dual_port_ram_0_douta_net_x0,
    ram_1_out => dual_port_ram_1_douta_net_x0,
    ram_2_out => dual_port_ram_2_douta_net_x0,
    ram_3_out => dual_port_ram_3_douta_net_x0,
    ram_4_out => dual_port_ram_4_douta_net_x0,
    valid => convert_to_bool_dout_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_a598ef7898 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
end structural;
-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH_struct
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_struct is
  port (
    data_enable_18_bit : in std_logic_vector( 1-1 downto 0 );
    data_in_18_bit : in std_logic_vector( 18-1 downto 0 );
    data_input_12_bit : in std_logic_vector( 12-1 downto 0 );
    write_enable_12_bit : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    kernel_line_gateway_conversion : out std_logic_vector( 12-1 downto 0 );
    kernel_output_gateway_conversion : out std_logic_vector( 128-1 downto 0 );
    kernel_serial_position_gateway_conversion : out std_logic_vector( 12-1 downto 0 );
    valid_kernel_output_gateway_conversion : out std_logic_vector( 1-1 downto 0 )
  );
end mh_struct;
architecture structural of mh_struct is 
  signal kernel_result_array_offset_op_net : std_logic_vector( 12-1 downto 0 );
  signal data_enable_18_bit_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_18_bit_net : std_logic_vector( 18-1 downto 0 );
  signal write_enable_12_bit_net : std_logic_vector( 1-1 downto 0 );
  signal data_input_12_bit_net : std_logic_vector( 12-1 downto 0 );
  signal output_enable_y_net : std_logic_vector( 1-1 downto 0 );
  signal output_or_block_y_net : std_logic_vector( 128-1 downto 0 );
  signal clk_net : std_logic;
  signal kernel_result_array_offset1_op_net : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal x12_bit_bin_value_6_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x5 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x8 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x4 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal data_valid_out_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_2_douta_net : std_logic_vector( 72-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_4_douta_net : std_logic_vector( 72-1 downto 0 );
  signal x12_bit_bin_value_4_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net : std_logic_vector( 18-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 72-1 downto 0 );
  signal x12_bit_bin_value_9_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net : std_logic_vector( 72-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_7_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_9_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_10_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_11_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_1_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_2_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_5_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_6_q_net : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_8_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal x12_bit_bin_value_3_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_2_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal convert_to_bool_dout_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_0_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_4_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
  signal dual_port_ram_3_douta_net_x0 : std_logic_vector( 72-1 downto 0 );
begin
  data_enable_18_bit_net <= data_enable_18_bit;
  data_in_18_bit_net <= data_in_18_bit;
  data_input_12_bit_net <= data_input_12_bit;
  kernel_line_gateway_conversion <= kernel_result_array_offset1_op_net;
  kernel_output_gateway_conversion <= output_or_block_y_net;
  kernel_serial_position_gateway_conversion <= kernel_result_array_offset_op_net;
  valid_kernel_output_gateway_conversion <= output_enable_y_net;
  write_enable_12_bit_net <= write_enable_12_bit;
  clk_net <= clk_1;
  ce_net <= ce_1;
  data_slicer : entity xil_defaultlib.mh_data_slicer 
  port map (
    data_in_ram_0 => dual_port_ram_0_douta_net,
    data_in_ram_1 => dual_port_ram_1_douta_net,
    data_in_ram_2 => dual_port_ram_2_douta_net,
    data_in_ram_3 => dual_port_ram_3_douta_net,
    data_in_ram_4 => dual_port_ram_4_douta_net,
    frame_valid_in => convert_to_bool_dout_net,
    kernel_data_in_ram_0 => dual_port_ram_0_douta_net_x0,
    kernel_data_in_ram_1 => dual_port_ram_1_douta_net_x0,
    kernel_data_in_ram_2 => dual_port_ram_2_douta_net_x0,
    kernel_data_in_ram_3 => dual_port_ram_3_douta_net_x0,
    kernel_data_in_ram_4 => dual_port_ram_4_douta_net_x0,
    kernel_valid_in => convert_to_bool_dout_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    frame_pixel_0_at_offset_0 => x12_bit_bin_value_0_q_net_x8,
    frame_pixel_1_at_offset_0 => x12_bit_bin_value_1_q_net_x7,
    frame_pixel_2_at_offset_0 => x12_bit_bin_value_2_q_net_x8,
    frame_pixel_3_at_offset_0 => x12_bit_bin_value_3_q_net_x8,
    frame_pixel_4_at_offset_0 => x12_bit_bin_value_4_q_net_x8,
    frame_pixel_5_at_offset_0 => x12_bit_bin_value_5_q_net_x8,
    frame_pixel_6_at_offset_0 => x12_bit_bin_value_6_q_net_x8,
    frame_pixel_7_at_offset_0 => x12_bit_bin_value_7_q_net_x8,
    frame_pixel_8_at_offset_0 => x12_bit_bin_value_8_q_net_x8,
    frame_pixel_9_at_offset_0 => x12_bit_bin_value_9_q_net_x8,
    frame_pixel_10_at_offset_0 => x12_bit_bin_value_10_q_net_x8,
    frame_pixel_11_at_offset_0 => x12_bit_bin_value_11_q_net_x8,
    frame_pixel_0_at_offset_1 => x12_bit_bin_value_0_q_net_x7,
    frame_pixel_1_at_offset_1 => x12_bit_bin_value_1_q_net_x8,
    frame_pixel_2_at_offset_1 => x12_bit_bin_value_2_q_net_x7,
    frame_pixel_3_at_offset_1 => x12_bit_bin_value_3_q_net_x7,
    frame_pixel_4_at_offset_1 => x12_bit_bin_value_4_q_net_x7,
    frame_pixel_5_at_offset_1 => x12_bit_bin_value_5_q_net_x7,
    frame_pixel_6_at_offset_1 => x12_bit_bin_value_6_q_net_x7,
    frame_pixel_7_at_offset_1 => x12_bit_bin_value_7_q_net_x6,
    frame_pixel_8_at_offset_1 => x12_bit_bin_value_8_q_net_x7,
    frame_pixel_9_at_offset_1 => x12_bit_bin_value_9_q_net_x7,
    frame_pixel_10_at_offset_1 => x12_bit_bin_value_10_q_net_x7,
    frame_pixel_11_at_offset_1 => x12_bit_bin_value_11_q_net_x7,
    frame_pixel_0_at_offset_2 => x12_bit_bin_value_0_q_net_x6,
    frame_pixel_1_at_offset_2 => x12_bit_bin_value_1_q_net_x6,
    frame_pixel_2_at_offset_2 => x12_bit_bin_value_2_q_net_x6,
    frame_pixel_3_at_offset_2 => x12_bit_bin_value_3_q_net_x6,
    frame_pixel_4_at_offset_2 => x12_bit_bin_value_4_q_net_x6,
    frame_pixel_5_at_offset_2 => x12_bit_bin_value_5_q_net_x6,
    frame_pixel_6_at_offset_2 => x12_bit_bin_value_6_q_net_x6,
    frame_pixel_7_at_offset_2 => x12_bit_bin_value_7_q_net_x7,
    frame_pixel_8_at_offset_2 => x12_bit_bin_value_8_q_net_x6,
    frame_pixel_9_at_offset_2 => x12_bit_bin_value_9_q_net_x6,
    frame_pixel_10_at_offset_2 => x12_bit_bin_value_10_q_net_x6,
    frame_pixel_11_at_offset_2 => x12_bit_bin_value_11_q_net_x6,
    frame_pixel_0_at_offset_3 => x12_bit_bin_value_0_q_net_x5,
    frame_pixel_1_at_offset_3 => x12_bit_bin_value_1_q_net_x5,
    frame_pixel_2_at_offset_3 => x12_bit_bin_value_2_q_net_x5,
    frame_pixel_3_at_offset_3 => x12_bit_bin_value_3_q_net_x5,
    frame_pixel_4_at_offset_3 => x12_bit_bin_value_4_q_net_x5,
    frame_pixel_5_at_offset_3 => x12_bit_bin_value_5_q_net_x5,
    frame_pixel_6_at_offset_3 => x12_bit_bin_value_6_q_net_x5,
    frame_pixel_7_at_offset_3 => x12_bit_bin_value_7_q_net_x5,
    frame_pixel_8_at_offset_3 => x12_bit_bin_value_8_q_net_x5,
    frame_pixel_9_at_offset_3 => x12_bit_bin_value_9_q_net_x5,
    frame_pixel_10_at_offset_3 => x12_bit_bin_value_10_q_net_x5,
    frame_pixel_11_at_offset_3 => x12_bit_bin_value_11_q_net_x5,
    frame_pixel_0_at_offset_4 => x12_bit_bin_value_0_q_net_x4,
    frame_pixel_1_at_offset_4 => x12_bit_bin_value_1_q_net_x4,
    frame_pixel_2_at_offset_4 => x12_bit_bin_value_2_q_net_x4,
    frame_pixel_3_at_offset_4 => x12_bit_bin_value_3_q_net_x4,
    frame_pixel_4_at_offset_4 => x12_bit_bin_value_4_q_net_x4,
    frame_pixel_5_at_offset_4 => x12_bit_bin_value_5_q_net_x4,
    frame_pixel_6_at_offset_4 => x12_bit_bin_value_6_q_net_x4,
    frame_pixel_7_at_offset_4 => x12_bit_bin_value_7_q_net_x4,
    frame_pixel_8_at_offset_4 => x12_bit_bin_value_8_q_net_x4,
    frame_pixel_9_at_offset_4 => x12_bit_bin_value_9_q_net_x4,
    frame_pixel_10_at_offset_4 => x12_bit_bin_value_10_q_net_x4,
    frame_pixel_11_at_offset_4 => x12_bit_bin_value_11_q_net_x4,
    weight_0_at_offset_0 => x12_bit_bin_value_0_q_net_x3,
    weight_1_at_offset_0 => x12_bit_bin_value_1_q_net_x3,
    weight_2_at_offset_0 => x12_bit_bin_value_2_q_net_x3,
    weight_3_at_offset_0 => x12_bit_bin_value_3_q_net_x3,
    weight_4_at_offset_0 => x12_bit_bin_value_4_q_net_x3,
    weight_5_at_offset_0 => x12_bit_bin_value_5_q_net_x3,
    weight_6_at_offset_0 => x12_bit_bin_value_6_q_net_x3,
    weight_7_at_offset_0 => x12_bit_bin_value_7_q_net_x3,
    weight_8_at_offset_0 => x12_bit_bin_value_8_q_net_x3,
    weight_9_at_offset_0 => x12_bit_bin_value_9_q_net_x3,
    weight_10_at_offset_0 => x12_bit_bin_value_10_q_net_x3,
    weight_11_at_offset_0 => x12_bit_bin_value_11_q_net_x3,
    weight_0_at_offset_1 => x12_bit_bin_value_0_q_net_x2,
    weight_1_at_offset_1 => x12_bit_bin_value_1_q_net_x2,
    weight_2_at_offset_1 => x12_bit_bin_value_2_q_net_x2,
    weight_3_at_offset_1 => x12_bit_bin_value_3_q_net_x2,
    weight_4_at_offset_1 => x12_bit_bin_value_4_q_net_x2,
    weight_5_at_offset_1 => x12_bit_bin_value_5_q_net_x2,
    weight_6_at_offset_1 => x12_bit_bin_value_6_q_net_x2,
    weight_7_at_offset_1 => x12_bit_bin_value_7_q_net_x2,
    weight_8_at_offset_1 => x12_bit_bin_value_8_q_net_x2,
    weight_9_at_offset_1 => x12_bit_bin_value_9_q_net_x2,
    weight_10_at_offset_1 => x12_bit_bin_value_10_q_net_x2,
    weight_11_at_offset_1 => x12_bit_bin_value_11_q_net_x2,
    weight_0_at_offset_2 => x12_bit_bin_value_0_q_net_x1,
    weight_1_at_offset_2 => x12_bit_bin_value_1_q_net_x1,
    weight_2_at_offset_2 => x12_bit_bin_value_2_q_net_x1,
    weight_3_at_offset_2 => x12_bit_bin_value_3_q_net_x1,
    weight_4_at_offset_2 => x12_bit_bin_value_4_q_net_x1,
    weight_5_at_offset_2 => x12_bit_bin_value_5_q_net_x1,
    weight_6_at_offset_2 => x12_bit_bin_value_6_q_net_x1,
    weight_7_at_offset_2 => x12_bit_bin_value_7_q_net_x1,
    weight_8_at_offset_2 => x12_bit_bin_value_8_q_net_x1,
    weight_9_at_offset_2 => x12_bit_bin_value_9_q_net_x1,
    weight_10_at_offset_2 => x12_bit_bin_value_10_q_net_x1,
    weight_11_at_offset_2 => x12_bit_bin_value_11_q_net_x1,
    weight_0_at_offset_3 => x12_bit_bin_value_0_q_net_x0,
    weight_1_at_offset_3 => x12_bit_bin_value_1_q_net_x0,
    weight_2_at_offset_3 => x12_bit_bin_value_2_q_net_x0,
    weight_3_at_offset_3 => x12_bit_bin_value_3_q_net_x0,
    weight_4_at_offset_3 => x12_bit_bin_value_4_q_net_x0,
    weight_5_at_offset_3 => x12_bit_bin_value_5_q_net_x0,
    weight_6_at_offset_3 => x12_bit_bin_value_6_q_net_x0,
    weight_7_at_offset_3 => x12_bit_bin_value_7_q_net_x0,
    weight_8_at_offset_3 => x12_bit_bin_value_8_q_net_x0,
    weight_9_at_offset_3 => x12_bit_bin_value_9_q_net_x0,
    weight_10_at_offset_3 => x12_bit_bin_value_10_q_net_x0,
    weight_11_at_offset_3 => x12_bit_bin_value_11_q_net_x0,
    weight_0_at_offset_4 => x12_bit_bin_value_0_q_net,
    weight_1_at_offset_4 => x12_bit_bin_value_1_q_net,
    weight_2_at_offset_4 => x12_bit_bin_value_2_q_net,
    weight_3_at_offset_4 => x12_bit_bin_value_3_q_net,
    weight_4_at_offset_4 => x12_bit_bin_value_4_q_net,
    weight_5_at_offset_4 => x12_bit_bin_value_5_q_net,
    weight_6_at_offset_4 => x12_bit_bin_value_6_q_net,
    weight_7_at_offset_4 => x12_bit_bin_value_7_q_net,
    weight_8_at_offset_4 => x12_bit_bin_value_8_q_net,
    weight_9_at_offset_4 => x12_bit_bin_value_9_q_net,
    weight_10_at_offset_4 => x12_bit_bin_value_10_q_net,
    weight_11_at_offset_4 => x12_bit_bin_value_11_q_net,
    valid_data => data_valid_out_delay_q_net
  );
  math : entity xil_defaultlib.mh_math 
  port map (
    in_pixel_0_at_offset_0 => x12_bit_bin_value_0_q_net_x8,
    in_pixel_1_at_offset_0 => x12_bit_bin_value_1_q_net_x7,
    in_pixel_2_at_offset_0 => x12_bit_bin_value_2_q_net_x8,
    in_pixel_3_at_offset_0 => x12_bit_bin_value_3_q_net_x8,
    in_pixel_4_at_offset_0 => x12_bit_bin_value_4_q_net_x8,
    in_pixel_5_at_offset_0 => x12_bit_bin_value_5_q_net_x8,
    in_pixel_6_at_offset_0 => x12_bit_bin_value_6_q_net_x8,
    in_pixel_7_at_offset_0 => x12_bit_bin_value_7_q_net_x8,
    in_pixel_8_at_offset_0 => x12_bit_bin_value_8_q_net_x8,
    in_pixel_9_at_offset_0 => x12_bit_bin_value_9_q_net_x8,
    in_pixel_10_at_offset_0 => x12_bit_bin_value_10_q_net_x8,
    in_pixel_11_at_offset_0 => x12_bit_bin_value_11_q_net_x8,
    in_pixel_0_at_offset_1 => x12_bit_bin_value_0_q_net_x7,
    in_pixel_1_at_offset_1 => x12_bit_bin_value_1_q_net_x8,
    in_pixel_2_at_offset_1 => x12_bit_bin_value_2_q_net_x7,
    in_pixel_3_at_offset_1 => x12_bit_bin_value_3_q_net_x7,
    in_pixel_4_at_offset_1 => x12_bit_bin_value_4_q_net_x7,
    in_pixel_5_at_offset_1 => x12_bit_bin_value_5_q_net_x7,
    in_pixel_6_at_offset_1 => x12_bit_bin_value_6_q_net_x7,
    in_pixel_7_at_offset_1 => x12_bit_bin_value_7_q_net_x6,
    in_pixel_8_at_offset_1 => x12_bit_bin_value_8_q_net_x7,
    in_pixel_9_at_offset_1 => x12_bit_bin_value_9_q_net_x7,
    in_pixel_10_at_offset_1 => x12_bit_bin_value_10_q_net_x7,
    in_pixel_11_at_offset_1 => x12_bit_bin_value_11_q_net_x7,
    in_pixel_0_at_offset_2 => x12_bit_bin_value_0_q_net_x6,
    in_pixel_1_at_offset_2 => x12_bit_bin_value_1_q_net_x6,
    in_pixel_2_at_offset_2 => x12_bit_bin_value_2_q_net_x6,
    in_pixel_3_at_offset_2 => x12_bit_bin_value_3_q_net_x6,
    in_pixel_4_at_offset_2 => x12_bit_bin_value_4_q_net_x6,
    in_pixel_5_at_offset_2 => x12_bit_bin_value_5_q_net_x6,
    in_pixel_6_at_offset_2 => x12_bit_bin_value_6_q_net_x6,
    in_pixel_7_at_offset_2 => x12_bit_bin_value_7_q_net_x7,
    in_pixel_8_at_offset_2 => x12_bit_bin_value_8_q_net_x6,
    in_pixel_9_at_offset_2 => x12_bit_bin_value_9_q_net_x6,
    in_pixel_10_at_offset_2 => x12_bit_bin_value_10_q_net_x6,
    in_pixel_11_at_offset_2 => x12_bit_bin_value_11_q_net_x6,
    in_pixel_0_at_offset_3 => x12_bit_bin_value_0_q_net_x5,
    in_pixel_1_at_offset_3 => x12_bit_bin_value_1_q_net_x5,
    in_pixel_2_at_offset_3 => x12_bit_bin_value_2_q_net_x5,
    in_pixel_3_at_offset_3 => x12_bit_bin_value_3_q_net_x5,
    in_pixel_4_at_offset_3 => x12_bit_bin_value_4_q_net_x5,
    in_pixel_5_at_offset_3 => x12_bit_bin_value_5_q_net_x5,
    in_pixel_6_at_offset_3 => x12_bit_bin_value_6_q_net_x5,
    in_pixel_7_at_offset_3 => x12_bit_bin_value_7_q_net_x5,
    in_pixel_8_at_offset_3 => x12_bit_bin_value_8_q_net_x5,
    in_pixel_9_at_offset_3 => x12_bit_bin_value_9_q_net_x5,
    in_pixel_10_at_offset_3 => x12_bit_bin_value_10_q_net_x5,
    in_pixel_11_at_offset_3 => x12_bit_bin_value_11_q_net_x5,
    in_pixel_0_at_offset_4 => x12_bit_bin_value_0_q_net_x4,
    in_pixel_1_at_offset_4 => x12_bit_bin_value_1_q_net_x4,
    in_pixel_2_at_offset_4 => x12_bit_bin_value_2_q_net_x4,
    in_pixel_3_at_offset_4 => x12_bit_bin_value_3_q_net_x4,
    in_pixel_4_at_offset_4 => x12_bit_bin_value_4_q_net_x4,
    in_pixel_5_at_offset_4 => x12_bit_bin_value_5_q_net_x4,
    in_pixel_6_at_offset_4 => x12_bit_bin_value_6_q_net_x4,
    in_pixel_7_at_offset_4 => x12_bit_bin_value_7_q_net_x4,
    in_pixel_8_at_offset_4 => x12_bit_bin_value_8_q_net_x4,
    in_pixel_9_at_offset_4 => x12_bit_bin_value_9_q_net_x4,
    in_pixel_10_at_offset_4 => x12_bit_bin_value_10_q_net_x4,
    in_pixel_11_at_offset_4 => x12_bit_bin_value_11_q_net_x4,
    in_weight_0_at_offset_0 => x12_bit_bin_value_0_q_net_x3,
    in_weight_1_at_offset_0 => x12_bit_bin_value_1_q_net_x3,
    in_weight_2_at_offset_0 => x12_bit_bin_value_2_q_net_x3,
    in_weight_3_at_offset_0 => x12_bit_bin_value_3_q_net_x3,
    in_weight_4_at_offset_0 => x12_bit_bin_value_4_q_net_x3,
    in_weight_5_at_offset_0 => x12_bit_bin_value_5_q_net_x3,
    in_weight_6_at_offset_0 => x12_bit_bin_value_6_q_net_x3,
    in_weight_7_at_offset_0 => x12_bit_bin_value_7_q_net_x3,
    in_weight_8_at_offset_0 => x12_bit_bin_value_8_q_net_x3,
    in_weight_9_at_offset_0 => x12_bit_bin_value_9_q_net_x3,
    in_weight_10_at_offset_0 => x12_bit_bin_value_10_q_net_x3,
    in_weight_11_at_offset_0 => x12_bit_bin_value_11_q_net_x3,
    in_weight_0_at_offset_1 => x12_bit_bin_value_0_q_net_x2,
    in_weight_1_at_offset_1 => x12_bit_bin_value_1_q_net_x2,
    in_weight_2_at_offset_1 => x12_bit_bin_value_2_q_net_x2,
    in_weight_3_at_offset_1 => x12_bit_bin_value_3_q_net_x2,
    in_weight_4_at_offset_1 => x12_bit_bin_value_4_q_net_x2,
    in_weight_5_at_offset_1 => x12_bit_bin_value_5_q_net_x2,
    in_weight_6_at_offset_1 => x12_bit_bin_value_6_q_net_x2,
    in_weight_7_at_offset_1 => x12_bit_bin_value_7_q_net_x2,
    in_weight_8_at_offset_1 => x12_bit_bin_value_8_q_net_x2,
    in_weight_9_at_offset_1 => x12_bit_bin_value_9_q_net_x2,
    in_weight_10_at_offset_1 => x12_bit_bin_value_10_q_net_x2,
    in_weight_11_at_offset_1 => x12_bit_bin_value_11_q_net_x2,
    in_weight_0_at_offset_2 => x12_bit_bin_value_0_q_net_x1,
    in_weight_1_at_offset_2 => x12_bit_bin_value_1_q_net_x1,
    in_weight_2_at_offset_2 => x12_bit_bin_value_2_q_net_x1,
    in_weight_3_at_offset_2 => x12_bit_bin_value_3_q_net_x1,
    in_weight_4_at_offset_2 => x12_bit_bin_value_4_q_net_x1,
    in_weight_5_at_offset_2 => x12_bit_bin_value_5_q_net_x1,
    in_weight_6_at_offset_2 => x12_bit_bin_value_6_q_net_x1,
    in_weight_7_at_offset_2 => x12_bit_bin_value_7_q_net_x1,
    in_weight_8_at_offset_2 => x12_bit_bin_value_8_q_net_x1,
    in_weight_9_at_offset_2 => x12_bit_bin_value_9_q_net_x1,
    in_weight_10_at_offset_2 => x12_bit_bin_value_10_q_net_x1,
    in_weight_11_at_offset_2 => x12_bit_bin_value_11_q_net_x1,
    in_weight_0_at_offset_3 => x12_bit_bin_value_0_q_net_x0,
    in_weight_1_at_offset_3 => x12_bit_bin_value_1_q_net_x0,
    in_weight_2_at_offset_3 => x12_bit_bin_value_2_q_net_x0,
    in_weight_3_at_offset_3 => x12_bit_bin_value_3_q_net_x0,
    in_weight_4_at_offset_3 => x12_bit_bin_value_4_q_net_x0,
    in_weight_5_at_offset_3 => x12_bit_bin_value_5_q_net_x0,
    in_weight_6_at_offset_3 => x12_bit_bin_value_6_q_net_x0,
    in_weight_7_at_offset_3 => x12_bit_bin_value_7_q_net_x0,
    in_weight_8_at_offset_3 => x12_bit_bin_value_8_q_net_x0,
    in_weight_9_at_offset_3 => x12_bit_bin_value_9_q_net_x0,
    in_weight_10_at_offset_3 => x12_bit_bin_value_10_q_net_x0,
    in_weight_11_at_offset_3 => x12_bit_bin_value_11_q_net_x0,
    in_weight_0_at_offset_4 => x12_bit_bin_value_0_q_net,
    in_weight_1_at_offset_4 => x12_bit_bin_value_1_q_net,
    in_weight_2_at_offset_4 => x12_bit_bin_value_2_q_net,
    in_weight_3_at_offset_4 => x12_bit_bin_value_3_q_net,
    in_weight_4_at_offset_4 => x12_bit_bin_value_4_q_net,
    in_weight_5_at_offset_4 => x12_bit_bin_value_5_q_net,
    in_weight_6_at_offset_4 => x12_bit_bin_value_6_q_net,
    in_weight_7_at_offset_4 => x12_bit_bin_value_7_q_net,
    in_weight_8_at_offset_4 => x12_bit_bin_value_8_q_net,
    in_weight_9_at_offset_4 => x12_bit_bin_value_9_q_net,
    in_weight_10_at_offset_4 => x12_bit_bin_value_10_q_net,
    in_weight_11_at_offset_4 => x12_bit_bin_value_11_q_net,
    valid_data_in => data_valid_out_delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    kernel_output => output_or_block_y_net,
    valid_kernel_output => output_enable_y_net,
    kernel_result_array_position => kernel_result_array_offset_op_net,
    kernel_result_row_depth_position => kernel_result_array_offset1_op_net
  );
  memory_manager : entity xil_defaultlib.mh_memory_manager 
  port map (
    x12_bit_spectrual_bin_in => data_input_12_bit_net,
    enable_in_spectrual => write_enable_12_bit_net,
    x18_bit_kernel_data_in => data_in_18_bit_net,
    enable_in_kernel => data_enable_18_bit_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    spectrual_ram_0_out => dual_port_ram_0_douta_net,
    spectrual_ram_1_out => dual_port_ram_1_douta_net,
    spectrual_ram_2_out => dual_port_ram_2_douta_net,
    spectrual_ram_3_out => dual_port_ram_3_douta_net,
    spectrual_ram_4_out => dual_port_ram_4_douta_net,
    spectrual_valid => convert_to_bool_dout_net,
    kernel_ram_0_out1 => dual_port_ram_0_douta_net_x0,
    kernel_ram_1_out1 => dual_port_ram_1_douta_net_x0,
    kernel_ram_2_out1 => dual_port_ram_2_douta_net_x0,
    kernel_ram_3_out1 => dual_port_ram_3_douta_net_x0,
    kernel_ram_4_out1 => dual_port_ram_4_douta_net_x0,
    kernel_valid => convert_to_bool_dout_net_x0
  );
end structural;
-- Generated from Simulink block 
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_default_clock_driver is
  port (
    mh_sysclk : in std_logic;
    mh_sysce : in std_logic;
    mh_sysclr : in std_logic;
    mh_clk1 : out std_logic;
    mh_ce1 : out std_logic
  );
end mh_default_clock_driver;
architecture structural of mh_default_clock_driver is 
begin
  clockdriver : entity xil_defaultlib.xlclockdriver 
  generic map (
    period => 1,
    log_2_period => 1
  )
  port map (
    sysclk => mh_sysclk,
    sysce => mh_sysce,
    sysclr => mh_sysclr,
    clk => mh_clk1,
    ce => mh_ce1
  );
end structural;
-- Generated from Simulink block 
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh is
  port (
    data_enable_18_bit : in std_logic;
    data_in_18_bit : in std_logic_vector( 18-1 downto 0 );
    data_input_12_bit : in std_logic_vector( 12-1 downto 0 );
    write_enable_12_bit : in std_logic;
    clk : in std_logic;
    kernel_line_gateway_conversion : out std_logic_vector( 12-1 downto 0 );
    kernel_output_gateway_conversion : out std_logic_vector( 128-1 downto 0 );
    kernel_serial_position_gateway_conversion : out std_logic_vector( 12-1 downto 0 );
    valid_kernel_output_gateway_conversion : out std_logic
  );
end mh;
architecture structural of mh is 
  attribute core_generation_info : string;
  attribute core_generation_info of structural : architecture is "mh,sysgen_core_2024_1,{,compilation=IP Catalog,block_icon_display=Default,family=zynquplus,part=xck26,speed=-2LV-c,package=sfvc784,synthesis_language=vhdl,hdl_library=xil_defaultlib,synthesis_strategy=Vivado Synthesis Defaults,implementation_strategy=Vivado Implementation Defaults,testbench=1,interface_doc=0,ce_clr=0,clock_period=10,system_simulink_period=1,waveform_viewer=1,axilite_interface=0,ip_catalog_plugin=0,hwcosim_burst_mode=0,simulation_time=10,accum=60,addsub=594,concat=2,constant=183,convert=7,counter=96,delay=2160,dpram=10,fifo=35,logical=312,mult=602,mux=184,relational=87,slice=172,}";
  signal clk_1_net : std_logic;
  signal ce_1_net : std_logic;
begin
  mh_default_clock_driver : entity xil_defaultlib.mh_default_clock_driver 
  port map (
    mh_sysclk => clk,
    mh_sysce => '1',
    mh_sysclr => '0',
    mh_clk1 => clk_1_net,
    mh_ce1 => ce_1_net
  );
  mh_struct : entity xil_defaultlib.mh_struct 
  port map (
    data_enable_18_bit(0) => data_enable_18_bit,
    data_in_18_bit => data_in_18_bit,
    data_input_12_bit => data_input_12_bit,
    write_enable_12_bit(0) => write_enable_12_bit,
    clk_1 => clk_1_net,
    ce_1 => ce_1_net,
    kernel_line_gateway_conversion => kernel_line_gateway_conversion,
    kernel_output_gateway_conversion => kernel_output_gateway_conversion,
    kernel_serial_position_gateway_conversion => kernel_serial_position_gateway_conversion,
    valid_kernel_output_gateway_conversion(0) => valid_kernel_output_gateway_conversion
  );
end structural;
