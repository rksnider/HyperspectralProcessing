-- Generated from Simulink block CMOS_Kernel_Memory_Sync/MH/Memory Manager/Kernel Memory Controller
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity mh_kernel_memory_controller is
  port (
    x18_bit_data_in : in std_logic_vector( 18-1 downto 0 );
    enable_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    data_out_72_bits : out std_logic_vector( 72-1 downto 0 );
    data_out_ready : out std_logic_vector( 1-1 downto 0 );
    data_address_out : out std_logic_vector( 9-1 downto 0 );
    ram_block_sel_out : out std_logic_vector( 3-1 downto 0 );
    memory_is_full : out std_logic_vector( 1-1 downto 0 )
  );
end mh_kernel_memory_controller;
architecture structural of mh_kernel_memory_controller is 
  signal ce_net : std_logic;
  signal multiple_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal final_add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal add_ram_sel_delay_1_q_net : std_logic_vector( 3-1 downto 0 );
  signal final_add_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal multiple_data_out_delay_q_net : std_logic_vector( 72-1 downto 0 );
  signal add_enable_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal data_in_18_bit_net : std_logic_vector( 18-1 downto 0 );
  signal data_points_per_line_op_net : std_logic_vector( 9-1 downto 0 );
  signal memory_full_delay_1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal data_out_delay_q_net : std_logic_vector( 9-1 downto 0 );
  signal add_line_delay_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal data_enable_18_bit_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_0_empty_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_3_empty_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_new_section_op_net : std_logic_vector( 1-1 downto 0 );
  signal check_new_line_delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_2_empty_net : std_logic_vector( 1-1 downto 0 );
  signal add_line_delay_1_q_net : std_logic_vector( 9-1 downto 0 );
  signal check_for_all_not_empty_y_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal offset_fifo_1_empty_net : std_logic_vector( 1-1 downto 0 );
  signal check_for_new_line_op_net : std_logic_vector( 1-1 downto 0 );
  signal add_ram_sel_delay_0_q_net : std_logic_vector( 3-1 downto 0 );
  signal and_for_new_section_y_net : std_logic_vector( 1-1 downto 0 );
  signal multiple_ram_sel_delay_q_net : std_logic_vector( 3-1 downto 0 );
  signal check_new_for_ands_q_net : std_logic_vector( 1-1 downto 0 );
  signal and_for_new_line_y_net : std_logic_vector( 1-1 downto 0 );
  signal compare_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 3-1 downto 0 );
  signal offset_fifo_0_dout_net : std_logic_vector( 18-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 1-1 downto 0 );
  signal check_if_full_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat_72_bit_packed_value_y_net : std_logic_vector( 72-1 downto 0 );
  signal mux_delay_enable_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 12-1 downto 0 );
  signal offset_fifo_3_dout_net : std_logic_vector( 18-1 downto 0 );
  signal offset_fifo_2_dout_net : std_logic_vector( 18-1 downto 0 );
  signal offset_fifo_1_dout_net : std_logic_vector( 18-1 downto 0 );
  signal ram_block_determination_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 9-1 downto 0 );
  signal convert_to_bool_dout_net : std_logic_vector( 1-1 downto 0 );
  signal convert_to_bool_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_2_op_net : std_logic_vector( 9-1 downto 0 );
  signal data_points_op_net : std_logic_vector( 9-1 downto 0 );
  signal write_enable_offset_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_compare_1_op_net : std_logic_vector( 9-1 downto 0 );
  signal convert_2_cycle_enable_to_1_cycle_op_net : std_logic_vector( 2-1 downto 0 );
  signal hold_up_read_out_op_net : std_logic_vector( 1-1 downto 0 );
  signal write_enable_offset_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal write_enable_offset_2_y_net : std_logic_vector( 1-1 downto 0 );
